magic
tech sky130A
magscale 1 2
timestamp 1750272439
<< checkpaint >>
rect -3932 -1804 16633 16492
<< viali >>
rect 1409 7837 1443 7871
rect 10977 7837 11011 7871
rect 1593 7701 1627 7735
rect 11161 7701 11195 7735
rect 6193 7497 6227 7531
rect 7205 7497 7239 7531
rect 1409 7361 1443 7395
rect 5825 7361 5859 7395
rect 6009 7361 6043 7395
rect 6561 7361 6595 7395
rect 7021 7361 7055 7395
rect 10977 7361 11011 7395
rect 6469 7293 6503 7327
rect 6929 7293 6963 7327
rect 1593 7225 1627 7259
rect 11161 7157 11195 7191
<< metal1 >>
rect 1104 12538 11592 12560
rect 1104 12486 2261 12538
rect 2313 12486 2325 12538
rect 2377 12486 2389 12538
rect 2441 12486 2453 12538
rect 2505 12486 2517 12538
rect 2569 12486 4883 12538
rect 4935 12486 4947 12538
rect 4999 12486 5011 12538
rect 5063 12486 5075 12538
rect 5127 12486 5139 12538
rect 5191 12486 7505 12538
rect 7557 12486 7569 12538
rect 7621 12486 7633 12538
rect 7685 12486 7697 12538
rect 7749 12486 7761 12538
rect 7813 12486 10127 12538
rect 10179 12486 10191 12538
rect 10243 12486 10255 12538
rect 10307 12486 10319 12538
rect 10371 12486 10383 12538
rect 10435 12486 11592 12538
rect 1104 12464 11592 12486
rect 1104 11994 11592 12016
rect 1104 11942 2921 11994
rect 2973 11942 2985 11994
rect 3037 11942 3049 11994
rect 3101 11942 3113 11994
rect 3165 11942 3177 11994
rect 3229 11942 5543 11994
rect 5595 11942 5607 11994
rect 5659 11942 5671 11994
rect 5723 11942 5735 11994
rect 5787 11942 5799 11994
rect 5851 11942 8165 11994
rect 8217 11942 8229 11994
rect 8281 11942 8293 11994
rect 8345 11942 8357 11994
rect 8409 11942 8421 11994
rect 8473 11942 10787 11994
rect 10839 11942 10851 11994
rect 10903 11942 10915 11994
rect 10967 11942 10979 11994
rect 11031 11942 11043 11994
rect 11095 11942 11592 11994
rect 1104 11920 11592 11942
rect 1104 11450 11592 11472
rect 1104 11398 2261 11450
rect 2313 11398 2325 11450
rect 2377 11398 2389 11450
rect 2441 11398 2453 11450
rect 2505 11398 2517 11450
rect 2569 11398 4883 11450
rect 4935 11398 4947 11450
rect 4999 11398 5011 11450
rect 5063 11398 5075 11450
rect 5127 11398 5139 11450
rect 5191 11398 7505 11450
rect 7557 11398 7569 11450
rect 7621 11398 7633 11450
rect 7685 11398 7697 11450
rect 7749 11398 7761 11450
rect 7813 11398 10127 11450
rect 10179 11398 10191 11450
rect 10243 11398 10255 11450
rect 10307 11398 10319 11450
rect 10371 11398 10383 11450
rect 10435 11398 11592 11450
rect 1104 11376 11592 11398
rect 1104 10906 11592 10928
rect 1104 10854 2921 10906
rect 2973 10854 2985 10906
rect 3037 10854 3049 10906
rect 3101 10854 3113 10906
rect 3165 10854 3177 10906
rect 3229 10854 5543 10906
rect 5595 10854 5607 10906
rect 5659 10854 5671 10906
rect 5723 10854 5735 10906
rect 5787 10854 5799 10906
rect 5851 10854 8165 10906
rect 8217 10854 8229 10906
rect 8281 10854 8293 10906
rect 8345 10854 8357 10906
rect 8409 10854 8421 10906
rect 8473 10854 10787 10906
rect 10839 10854 10851 10906
rect 10903 10854 10915 10906
rect 10967 10854 10979 10906
rect 11031 10854 11043 10906
rect 11095 10854 11592 10906
rect 1104 10832 11592 10854
rect 1104 10362 11592 10384
rect 1104 10310 2261 10362
rect 2313 10310 2325 10362
rect 2377 10310 2389 10362
rect 2441 10310 2453 10362
rect 2505 10310 2517 10362
rect 2569 10310 4883 10362
rect 4935 10310 4947 10362
rect 4999 10310 5011 10362
rect 5063 10310 5075 10362
rect 5127 10310 5139 10362
rect 5191 10310 7505 10362
rect 7557 10310 7569 10362
rect 7621 10310 7633 10362
rect 7685 10310 7697 10362
rect 7749 10310 7761 10362
rect 7813 10310 10127 10362
rect 10179 10310 10191 10362
rect 10243 10310 10255 10362
rect 10307 10310 10319 10362
rect 10371 10310 10383 10362
rect 10435 10310 11592 10362
rect 1104 10288 11592 10310
rect 1104 9818 11592 9840
rect 1104 9766 2921 9818
rect 2973 9766 2985 9818
rect 3037 9766 3049 9818
rect 3101 9766 3113 9818
rect 3165 9766 3177 9818
rect 3229 9766 5543 9818
rect 5595 9766 5607 9818
rect 5659 9766 5671 9818
rect 5723 9766 5735 9818
rect 5787 9766 5799 9818
rect 5851 9766 8165 9818
rect 8217 9766 8229 9818
rect 8281 9766 8293 9818
rect 8345 9766 8357 9818
rect 8409 9766 8421 9818
rect 8473 9766 10787 9818
rect 10839 9766 10851 9818
rect 10903 9766 10915 9818
rect 10967 9766 10979 9818
rect 11031 9766 11043 9818
rect 11095 9766 11592 9818
rect 1104 9744 11592 9766
rect 1104 9274 11592 9296
rect 1104 9222 2261 9274
rect 2313 9222 2325 9274
rect 2377 9222 2389 9274
rect 2441 9222 2453 9274
rect 2505 9222 2517 9274
rect 2569 9222 4883 9274
rect 4935 9222 4947 9274
rect 4999 9222 5011 9274
rect 5063 9222 5075 9274
rect 5127 9222 5139 9274
rect 5191 9222 7505 9274
rect 7557 9222 7569 9274
rect 7621 9222 7633 9274
rect 7685 9222 7697 9274
rect 7749 9222 7761 9274
rect 7813 9222 10127 9274
rect 10179 9222 10191 9274
rect 10243 9222 10255 9274
rect 10307 9222 10319 9274
rect 10371 9222 10383 9274
rect 10435 9222 11592 9274
rect 1104 9200 11592 9222
rect 1104 8730 11592 8752
rect 1104 8678 2921 8730
rect 2973 8678 2985 8730
rect 3037 8678 3049 8730
rect 3101 8678 3113 8730
rect 3165 8678 3177 8730
rect 3229 8678 5543 8730
rect 5595 8678 5607 8730
rect 5659 8678 5671 8730
rect 5723 8678 5735 8730
rect 5787 8678 5799 8730
rect 5851 8678 8165 8730
rect 8217 8678 8229 8730
rect 8281 8678 8293 8730
rect 8345 8678 8357 8730
rect 8409 8678 8421 8730
rect 8473 8678 10787 8730
rect 10839 8678 10851 8730
rect 10903 8678 10915 8730
rect 10967 8678 10979 8730
rect 11031 8678 11043 8730
rect 11095 8678 11592 8730
rect 1104 8656 11592 8678
rect 1104 8186 11592 8208
rect 1104 8134 2261 8186
rect 2313 8134 2325 8186
rect 2377 8134 2389 8186
rect 2441 8134 2453 8186
rect 2505 8134 2517 8186
rect 2569 8134 4883 8186
rect 4935 8134 4947 8186
rect 4999 8134 5011 8186
rect 5063 8134 5075 8186
rect 5127 8134 5139 8186
rect 5191 8134 7505 8186
rect 7557 8134 7569 8186
rect 7621 8134 7633 8186
rect 7685 8134 7697 8186
rect 7749 8134 7761 8186
rect 7813 8134 10127 8186
rect 10179 8134 10191 8186
rect 10243 8134 10255 8186
rect 10307 8134 10319 8186
rect 10371 8134 10383 8186
rect 10435 8134 11592 8186
rect 1104 8112 11592 8134
rect 842 7828 848 7880
rect 900 7868 906 7880
rect 1397 7871 1455 7877
rect 1397 7868 1409 7871
rect 900 7840 1409 7868
rect 900 7828 906 7840
rect 1397 7837 1409 7840
rect 1443 7837 1455 7871
rect 1397 7831 1455 7837
rect 7190 7828 7196 7880
rect 7248 7868 7254 7880
rect 10965 7871 11023 7877
rect 10965 7868 10977 7871
rect 7248 7840 10977 7868
rect 7248 7828 7254 7840
rect 10965 7837 10977 7840
rect 11011 7837 11023 7871
rect 10965 7831 11023 7837
rect 1578 7692 1584 7744
rect 1636 7692 1642 7744
rect 11149 7735 11207 7741
rect 11149 7701 11161 7735
rect 11195 7732 11207 7735
rect 11238 7732 11244 7744
rect 11195 7704 11244 7732
rect 11195 7701 11207 7704
rect 11149 7695 11207 7701
rect 11238 7692 11244 7704
rect 11296 7692 11302 7744
rect 1104 7642 11592 7664
rect 1104 7590 2921 7642
rect 2973 7590 2985 7642
rect 3037 7590 3049 7642
rect 3101 7590 3113 7642
rect 3165 7590 3177 7642
rect 3229 7590 5543 7642
rect 5595 7590 5607 7642
rect 5659 7590 5671 7642
rect 5723 7590 5735 7642
rect 5787 7590 5799 7642
rect 5851 7590 8165 7642
rect 8217 7590 8229 7642
rect 8281 7590 8293 7642
rect 8345 7590 8357 7642
rect 8409 7590 8421 7642
rect 8473 7590 10787 7642
rect 10839 7590 10851 7642
rect 10903 7590 10915 7642
rect 10967 7590 10979 7642
rect 11031 7590 11043 7642
rect 11095 7590 11592 7642
rect 1104 7568 11592 7590
rect 6181 7531 6239 7537
rect 6181 7497 6193 7531
rect 6227 7528 6239 7531
rect 6227 7500 6914 7528
rect 6227 7497 6239 7500
rect 6181 7491 6239 7497
rect 5828 7432 6592 7460
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1578 7352 1584 7404
rect 1636 7392 1642 7404
rect 5828 7401 5856 7432
rect 6564 7401 6592 7432
rect 5813 7395 5871 7401
rect 5813 7392 5825 7395
rect 1636 7364 5825 7392
rect 1636 7352 1642 7364
rect 5813 7361 5825 7364
rect 5859 7361 5871 7395
rect 5813 7355 5871 7361
rect 5997 7395 6055 7401
rect 5997 7361 6009 7395
rect 6043 7361 6055 7395
rect 5997 7355 6055 7361
rect 6549 7395 6607 7401
rect 6549 7361 6561 7395
rect 6595 7361 6607 7395
rect 6886 7392 6914 7500
rect 7190 7488 7196 7540
rect 7248 7488 7254 7540
rect 7009 7395 7067 7401
rect 7009 7392 7021 7395
rect 6886 7364 7021 7392
rect 6549 7355 6607 7361
rect 7009 7361 7021 7364
rect 7055 7361 7067 7395
rect 7009 7355 7067 7361
rect 10965 7395 11023 7401
rect 10965 7361 10977 7395
rect 11011 7361 11023 7395
rect 10965 7355 11023 7361
rect 6012 7324 6040 7355
rect 6457 7327 6515 7333
rect 6457 7324 6469 7327
rect 1596 7296 6469 7324
rect 1596 7265 1624 7296
rect 6457 7293 6469 7296
rect 6503 7293 6515 7327
rect 6457 7287 6515 7293
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7324 6975 7327
rect 10980 7324 11008 7355
rect 6963 7296 11008 7324
rect 6963 7293 6975 7296
rect 6917 7287 6975 7293
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7225 1639 7259
rect 1581 7219 1639 7225
rect 11146 7148 11152 7200
rect 11204 7148 11210 7200
rect 1104 7098 11592 7120
rect 1104 7046 2261 7098
rect 2313 7046 2325 7098
rect 2377 7046 2389 7098
rect 2441 7046 2453 7098
rect 2505 7046 2517 7098
rect 2569 7046 4883 7098
rect 4935 7046 4947 7098
rect 4999 7046 5011 7098
rect 5063 7046 5075 7098
rect 5127 7046 5139 7098
rect 5191 7046 7505 7098
rect 7557 7046 7569 7098
rect 7621 7046 7633 7098
rect 7685 7046 7697 7098
rect 7749 7046 7761 7098
rect 7813 7046 10127 7098
rect 10179 7046 10191 7098
rect 10243 7046 10255 7098
rect 10307 7046 10319 7098
rect 10371 7046 10383 7098
rect 10435 7046 11592 7098
rect 1104 7024 11592 7046
rect 1104 6554 11592 6576
rect 1104 6502 2921 6554
rect 2973 6502 2985 6554
rect 3037 6502 3049 6554
rect 3101 6502 3113 6554
rect 3165 6502 3177 6554
rect 3229 6502 5543 6554
rect 5595 6502 5607 6554
rect 5659 6502 5671 6554
rect 5723 6502 5735 6554
rect 5787 6502 5799 6554
rect 5851 6502 8165 6554
rect 8217 6502 8229 6554
rect 8281 6502 8293 6554
rect 8345 6502 8357 6554
rect 8409 6502 8421 6554
rect 8473 6502 10787 6554
rect 10839 6502 10851 6554
rect 10903 6502 10915 6554
rect 10967 6502 10979 6554
rect 11031 6502 11043 6554
rect 11095 6502 11592 6554
rect 1104 6480 11592 6502
rect 1104 6010 11592 6032
rect 1104 5958 2261 6010
rect 2313 5958 2325 6010
rect 2377 5958 2389 6010
rect 2441 5958 2453 6010
rect 2505 5958 2517 6010
rect 2569 5958 4883 6010
rect 4935 5958 4947 6010
rect 4999 5958 5011 6010
rect 5063 5958 5075 6010
rect 5127 5958 5139 6010
rect 5191 5958 7505 6010
rect 7557 5958 7569 6010
rect 7621 5958 7633 6010
rect 7685 5958 7697 6010
rect 7749 5958 7761 6010
rect 7813 5958 10127 6010
rect 10179 5958 10191 6010
rect 10243 5958 10255 6010
rect 10307 5958 10319 6010
rect 10371 5958 10383 6010
rect 10435 5958 11592 6010
rect 1104 5936 11592 5958
rect 1104 5466 11592 5488
rect 1104 5414 2921 5466
rect 2973 5414 2985 5466
rect 3037 5414 3049 5466
rect 3101 5414 3113 5466
rect 3165 5414 3177 5466
rect 3229 5414 5543 5466
rect 5595 5414 5607 5466
rect 5659 5414 5671 5466
rect 5723 5414 5735 5466
rect 5787 5414 5799 5466
rect 5851 5414 8165 5466
rect 8217 5414 8229 5466
rect 8281 5414 8293 5466
rect 8345 5414 8357 5466
rect 8409 5414 8421 5466
rect 8473 5414 10787 5466
rect 10839 5414 10851 5466
rect 10903 5414 10915 5466
rect 10967 5414 10979 5466
rect 11031 5414 11043 5466
rect 11095 5414 11592 5466
rect 1104 5392 11592 5414
rect 1104 4922 11592 4944
rect 1104 4870 2261 4922
rect 2313 4870 2325 4922
rect 2377 4870 2389 4922
rect 2441 4870 2453 4922
rect 2505 4870 2517 4922
rect 2569 4870 4883 4922
rect 4935 4870 4947 4922
rect 4999 4870 5011 4922
rect 5063 4870 5075 4922
rect 5127 4870 5139 4922
rect 5191 4870 7505 4922
rect 7557 4870 7569 4922
rect 7621 4870 7633 4922
rect 7685 4870 7697 4922
rect 7749 4870 7761 4922
rect 7813 4870 10127 4922
rect 10179 4870 10191 4922
rect 10243 4870 10255 4922
rect 10307 4870 10319 4922
rect 10371 4870 10383 4922
rect 10435 4870 11592 4922
rect 1104 4848 11592 4870
rect 1104 4378 11592 4400
rect 1104 4326 2921 4378
rect 2973 4326 2985 4378
rect 3037 4326 3049 4378
rect 3101 4326 3113 4378
rect 3165 4326 3177 4378
rect 3229 4326 5543 4378
rect 5595 4326 5607 4378
rect 5659 4326 5671 4378
rect 5723 4326 5735 4378
rect 5787 4326 5799 4378
rect 5851 4326 8165 4378
rect 8217 4326 8229 4378
rect 8281 4326 8293 4378
rect 8345 4326 8357 4378
rect 8409 4326 8421 4378
rect 8473 4326 10787 4378
rect 10839 4326 10851 4378
rect 10903 4326 10915 4378
rect 10967 4326 10979 4378
rect 11031 4326 11043 4378
rect 11095 4326 11592 4378
rect 1104 4304 11592 4326
rect 1104 3834 11592 3856
rect 1104 3782 2261 3834
rect 2313 3782 2325 3834
rect 2377 3782 2389 3834
rect 2441 3782 2453 3834
rect 2505 3782 2517 3834
rect 2569 3782 4883 3834
rect 4935 3782 4947 3834
rect 4999 3782 5011 3834
rect 5063 3782 5075 3834
rect 5127 3782 5139 3834
rect 5191 3782 7505 3834
rect 7557 3782 7569 3834
rect 7621 3782 7633 3834
rect 7685 3782 7697 3834
rect 7749 3782 7761 3834
rect 7813 3782 10127 3834
rect 10179 3782 10191 3834
rect 10243 3782 10255 3834
rect 10307 3782 10319 3834
rect 10371 3782 10383 3834
rect 10435 3782 11592 3834
rect 1104 3760 11592 3782
rect 1104 3290 11592 3312
rect 1104 3238 2921 3290
rect 2973 3238 2985 3290
rect 3037 3238 3049 3290
rect 3101 3238 3113 3290
rect 3165 3238 3177 3290
rect 3229 3238 5543 3290
rect 5595 3238 5607 3290
rect 5659 3238 5671 3290
rect 5723 3238 5735 3290
rect 5787 3238 5799 3290
rect 5851 3238 8165 3290
rect 8217 3238 8229 3290
rect 8281 3238 8293 3290
rect 8345 3238 8357 3290
rect 8409 3238 8421 3290
rect 8473 3238 10787 3290
rect 10839 3238 10851 3290
rect 10903 3238 10915 3290
rect 10967 3238 10979 3290
rect 11031 3238 11043 3290
rect 11095 3238 11592 3290
rect 1104 3216 11592 3238
rect 1104 2746 11592 2768
rect 1104 2694 2261 2746
rect 2313 2694 2325 2746
rect 2377 2694 2389 2746
rect 2441 2694 2453 2746
rect 2505 2694 2517 2746
rect 2569 2694 4883 2746
rect 4935 2694 4947 2746
rect 4999 2694 5011 2746
rect 5063 2694 5075 2746
rect 5127 2694 5139 2746
rect 5191 2694 7505 2746
rect 7557 2694 7569 2746
rect 7621 2694 7633 2746
rect 7685 2694 7697 2746
rect 7749 2694 7761 2746
rect 7813 2694 10127 2746
rect 10179 2694 10191 2746
rect 10243 2694 10255 2746
rect 10307 2694 10319 2746
rect 10371 2694 10383 2746
rect 10435 2694 11592 2746
rect 1104 2672 11592 2694
rect 1104 2202 11592 2224
rect 1104 2150 2921 2202
rect 2973 2150 2985 2202
rect 3037 2150 3049 2202
rect 3101 2150 3113 2202
rect 3165 2150 3177 2202
rect 3229 2150 5543 2202
rect 5595 2150 5607 2202
rect 5659 2150 5671 2202
rect 5723 2150 5735 2202
rect 5787 2150 5799 2202
rect 5851 2150 8165 2202
rect 8217 2150 8229 2202
rect 8281 2150 8293 2202
rect 8345 2150 8357 2202
rect 8409 2150 8421 2202
rect 8473 2150 10787 2202
rect 10839 2150 10851 2202
rect 10903 2150 10915 2202
rect 10967 2150 10979 2202
rect 11031 2150 11043 2202
rect 11095 2150 11592 2202
rect 1104 2128 11592 2150
<< via1 >>
rect 2261 12486 2313 12538
rect 2325 12486 2377 12538
rect 2389 12486 2441 12538
rect 2453 12486 2505 12538
rect 2517 12486 2569 12538
rect 4883 12486 4935 12538
rect 4947 12486 4999 12538
rect 5011 12486 5063 12538
rect 5075 12486 5127 12538
rect 5139 12486 5191 12538
rect 7505 12486 7557 12538
rect 7569 12486 7621 12538
rect 7633 12486 7685 12538
rect 7697 12486 7749 12538
rect 7761 12486 7813 12538
rect 10127 12486 10179 12538
rect 10191 12486 10243 12538
rect 10255 12486 10307 12538
rect 10319 12486 10371 12538
rect 10383 12486 10435 12538
rect 2921 11942 2973 11994
rect 2985 11942 3037 11994
rect 3049 11942 3101 11994
rect 3113 11942 3165 11994
rect 3177 11942 3229 11994
rect 5543 11942 5595 11994
rect 5607 11942 5659 11994
rect 5671 11942 5723 11994
rect 5735 11942 5787 11994
rect 5799 11942 5851 11994
rect 8165 11942 8217 11994
rect 8229 11942 8281 11994
rect 8293 11942 8345 11994
rect 8357 11942 8409 11994
rect 8421 11942 8473 11994
rect 10787 11942 10839 11994
rect 10851 11942 10903 11994
rect 10915 11942 10967 11994
rect 10979 11942 11031 11994
rect 11043 11942 11095 11994
rect 2261 11398 2313 11450
rect 2325 11398 2377 11450
rect 2389 11398 2441 11450
rect 2453 11398 2505 11450
rect 2517 11398 2569 11450
rect 4883 11398 4935 11450
rect 4947 11398 4999 11450
rect 5011 11398 5063 11450
rect 5075 11398 5127 11450
rect 5139 11398 5191 11450
rect 7505 11398 7557 11450
rect 7569 11398 7621 11450
rect 7633 11398 7685 11450
rect 7697 11398 7749 11450
rect 7761 11398 7813 11450
rect 10127 11398 10179 11450
rect 10191 11398 10243 11450
rect 10255 11398 10307 11450
rect 10319 11398 10371 11450
rect 10383 11398 10435 11450
rect 2921 10854 2973 10906
rect 2985 10854 3037 10906
rect 3049 10854 3101 10906
rect 3113 10854 3165 10906
rect 3177 10854 3229 10906
rect 5543 10854 5595 10906
rect 5607 10854 5659 10906
rect 5671 10854 5723 10906
rect 5735 10854 5787 10906
rect 5799 10854 5851 10906
rect 8165 10854 8217 10906
rect 8229 10854 8281 10906
rect 8293 10854 8345 10906
rect 8357 10854 8409 10906
rect 8421 10854 8473 10906
rect 10787 10854 10839 10906
rect 10851 10854 10903 10906
rect 10915 10854 10967 10906
rect 10979 10854 11031 10906
rect 11043 10854 11095 10906
rect 2261 10310 2313 10362
rect 2325 10310 2377 10362
rect 2389 10310 2441 10362
rect 2453 10310 2505 10362
rect 2517 10310 2569 10362
rect 4883 10310 4935 10362
rect 4947 10310 4999 10362
rect 5011 10310 5063 10362
rect 5075 10310 5127 10362
rect 5139 10310 5191 10362
rect 7505 10310 7557 10362
rect 7569 10310 7621 10362
rect 7633 10310 7685 10362
rect 7697 10310 7749 10362
rect 7761 10310 7813 10362
rect 10127 10310 10179 10362
rect 10191 10310 10243 10362
rect 10255 10310 10307 10362
rect 10319 10310 10371 10362
rect 10383 10310 10435 10362
rect 2921 9766 2973 9818
rect 2985 9766 3037 9818
rect 3049 9766 3101 9818
rect 3113 9766 3165 9818
rect 3177 9766 3229 9818
rect 5543 9766 5595 9818
rect 5607 9766 5659 9818
rect 5671 9766 5723 9818
rect 5735 9766 5787 9818
rect 5799 9766 5851 9818
rect 8165 9766 8217 9818
rect 8229 9766 8281 9818
rect 8293 9766 8345 9818
rect 8357 9766 8409 9818
rect 8421 9766 8473 9818
rect 10787 9766 10839 9818
rect 10851 9766 10903 9818
rect 10915 9766 10967 9818
rect 10979 9766 11031 9818
rect 11043 9766 11095 9818
rect 2261 9222 2313 9274
rect 2325 9222 2377 9274
rect 2389 9222 2441 9274
rect 2453 9222 2505 9274
rect 2517 9222 2569 9274
rect 4883 9222 4935 9274
rect 4947 9222 4999 9274
rect 5011 9222 5063 9274
rect 5075 9222 5127 9274
rect 5139 9222 5191 9274
rect 7505 9222 7557 9274
rect 7569 9222 7621 9274
rect 7633 9222 7685 9274
rect 7697 9222 7749 9274
rect 7761 9222 7813 9274
rect 10127 9222 10179 9274
rect 10191 9222 10243 9274
rect 10255 9222 10307 9274
rect 10319 9222 10371 9274
rect 10383 9222 10435 9274
rect 2921 8678 2973 8730
rect 2985 8678 3037 8730
rect 3049 8678 3101 8730
rect 3113 8678 3165 8730
rect 3177 8678 3229 8730
rect 5543 8678 5595 8730
rect 5607 8678 5659 8730
rect 5671 8678 5723 8730
rect 5735 8678 5787 8730
rect 5799 8678 5851 8730
rect 8165 8678 8217 8730
rect 8229 8678 8281 8730
rect 8293 8678 8345 8730
rect 8357 8678 8409 8730
rect 8421 8678 8473 8730
rect 10787 8678 10839 8730
rect 10851 8678 10903 8730
rect 10915 8678 10967 8730
rect 10979 8678 11031 8730
rect 11043 8678 11095 8730
rect 2261 8134 2313 8186
rect 2325 8134 2377 8186
rect 2389 8134 2441 8186
rect 2453 8134 2505 8186
rect 2517 8134 2569 8186
rect 4883 8134 4935 8186
rect 4947 8134 4999 8186
rect 5011 8134 5063 8186
rect 5075 8134 5127 8186
rect 5139 8134 5191 8186
rect 7505 8134 7557 8186
rect 7569 8134 7621 8186
rect 7633 8134 7685 8186
rect 7697 8134 7749 8186
rect 7761 8134 7813 8186
rect 10127 8134 10179 8186
rect 10191 8134 10243 8186
rect 10255 8134 10307 8186
rect 10319 8134 10371 8186
rect 10383 8134 10435 8186
rect 848 7828 900 7880
rect 7196 7828 7248 7880
rect 1584 7735 1636 7744
rect 1584 7701 1593 7735
rect 1593 7701 1627 7735
rect 1627 7701 1636 7735
rect 1584 7692 1636 7701
rect 11244 7692 11296 7744
rect 2921 7590 2973 7642
rect 2985 7590 3037 7642
rect 3049 7590 3101 7642
rect 3113 7590 3165 7642
rect 3177 7590 3229 7642
rect 5543 7590 5595 7642
rect 5607 7590 5659 7642
rect 5671 7590 5723 7642
rect 5735 7590 5787 7642
rect 5799 7590 5851 7642
rect 8165 7590 8217 7642
rect 8229 7590 8281 7642
rect 8293 7590 8345 7642
rect 8357 7590 8409 7642
rect 8421 7590 8473 7642
rect 10787 7590 10839 7642
rect 10851 7590 10903 7642
rect 10915 7590 10967 7642
rect 10979 7590 11031 7642
rect 11043 7590 11095 7642
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1584 7352 1636 7404
rect 7196 7531 7248 7540
rect 7196 7497 7205 7531
rect 7205 7497 7239 7531
rect 7239 7497 7248 7531
rect 7196 7488 7248 7497
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 2261 7046 2313 7098
rect 2325 7046 2377 7098
rect 2389 7046 2441 7098
rect 2453 7046 2505 7098
rect 2517 7046 2569 7098
rect 4883 7046 4935 7098
rect 4947 7046 4999 7098
rect 5011 7046 5063 7098
rect 5075 7046 5127 7098
rect 5139 7046 5191 7098
rect 7505 7046 7557 7098
rect 7569 7046 7621 7098
rect 7633 7046 7685 7098
rect 7697 7046 7749 7098
rect 7761 7046 7813 7098
rect 10127 7046 10179 7098
rect 10191 7046 10243 7098
rect 10255 7046 10307 7098
rect 10319 7046 10371 7098
rect 10383 7046 10435 7098
rect 2921 6502 2973 6554
rect 2985 6502 3037 6554
rect 3049 6502 3101 6554
rect 3113 6502 3165 6554
rect 3177 6502 3229 6554
rect 5543 6502 5595 6554
rect 5607 6502 5659 6554
rect 5671 6502 5723 6554
rect 5735 6502 5787 6554
rect 5799 6502 5851 6554
rect 8165 6502 8217 6554
rect 8229 6502 8281 6554
rect 8293 6502 8345 6554
rect 8357 6502 8409 6554
rect 8421 6502 8473 6554
rect 10787 6502 10839 6554
rect 10851 6502 10903 6554
rect 10915 6502 10967 6554
rect 10979 6502 11031 6554
rect 11043 6502 11095 6554
rect 2261 5958 2313 6010
rect 2325 5958 2377 6010
rect 2389 5958 2441 6010
rect 2453 5958 2505 6010
rect 2517 5958 2569 6010
rect 4883 5958 4935 6010
rect 4947 5958 4999 6010
rect 5011 5958 5063 6010
rect 5075 5958 5127 6010
rect 5139 5958 5191 6010
rect 7505 5958 7557 6010
rect 7569 5958 7621 6010
rect 7633 5958 7685 6010
rect 7697 5958 7749 6010
rect 7761 5958 7813 6010
rect 10127 5958 10179 6010
rect 10191 5958 10243 6010
rect 10255 5958 10307 6010
rect 10319 5958 10371 6010
rect 10383 5958 10435 6010
rect 2921 5414 2973 5466
rect 2985 5414 3037 5466
rect 3049 5414 3101 5466
rect 3113 5414 3165 5466
rect 3177 5414 3229 5466
rect 5543 5414 5595 5466
rect 5607 5414 5659 5466
rect 5671 5414 5723 5466
rect 5735 5414 5787 5466
rect 5799 5414 5851 5466
rect 8165 5414 8217 5466
rect 8229 5414 8281 5466
rect 8293 5414 8345 5466
rect 8357 5414 8409 5466
rect 8421 5414 8473 5466
rect 10787 5414 10839 5466
rect 10851 5414 10903 5466
rect 10915 5414 10967 5466
rect 10979 5414 11031 5466
rect 11043 5414 11095 5466
rect 2261 4870 2313 4922
rect 2325 4870 2377 4922
rect 2389 4870 2441 4922
rect 2453 4870 2505 4922
rect 2517 4870 2569 4922
rect 4883 4870 4935 4922
rect 4947 4870 4999 4922
rect 5011 4870 5063 4922
rect 5075 4870 5127 4922
rect 5139 4870 5191 4922
rect 7505 4870 7557 4922
rect 7569 4870 7621 4922
rect 7633 4870 7685 4922
rect 7697 4870 7749 4922
rect 7761 4870 7813 4922
rect 10127 4870 10179 4922
rect 10191 4870 10243 4922
rect 10255 4870 10307 4922
rect 10319 4870 10371 4922
rect 10383 4870 10435 4922
rect 2921 4326 2973 4378
rect 2985 4326 3037 4378
rect 3049 4326 3101 4378
rect 3113 4326 3165 4378
rect 3177 4326 3229 4378
rect 5543 4326 5595 4378
rect 5607 4326 5659 4378
rect 5671 4326 5723 4378
rect 5735 4326 5787 4378
rect 5799 4326 5851 4378
rect 8165 4326 8217 4378
rect 8229 4326 8281 4378
rect 8293 4326 8345 4378
rect 8357 4326 8409 4378
rect 8421 4326 8473 4378
rect 10787 4326 10839 4378
rect 10851 4326 10903 4378
rect 10915 4326 10967 4378
rect 10979 4326 11031 4378
rect 11043 4326 11095 4378
rect 2261 3782 2313 3834
rect 2325 3782 2377 3834
rect 2389 3782 2441 3834
rect 2453 3782 2505 3834
rect 2517 3782 2569 3834
rect 4883 3782 4935 3834
rect 4947 3782 4999 3834
rect 5011 3782 5063 3834
rect 5075 3782 5127 3834
rect 5139 3782 5191 3834
rect 7505 3782 7557 3834
rect 7569 3782 7621 3834
rect 7633 3782 7685 3834
rect 7697 3782 7749 3834
rect 7761 3782 7813 3834
rect 10127 3782 10179 3834
rect 10191 3782 10243 3834
rect 10255 3782 10307 3834
rect 10319 3782 10371 3834
rect 10383 3782 10435 3834
rect 2921 3238 2973 3290
rect 2985 3238 3037 3290
rect 3049 3238 3101 3290
rect 3113 3238 3165 3290
rect 3177 3238 3229 3290
rect 5543 3238 5595 3290
rect 5607 3238 5659 3290
rect 5671 3238 5723 3290
rect 5735 3238 5787 3290
rect 5799 3238 5851 3290
rect 8165 3238 8217 3290
rect 8229 3238 8281 3290
rect 8293 3238 8345 3290
rect 8357 3238 8409 3290
rect 8421 3238 8473 3290
rect 10787 3238 10839 3290
rect 10851 3238 10903 3290
rect 10915 3238 10967 3290
rect 10979 3238 11031 3290
rect 11043 3238 11095 3290
rect 2261 2694 2313 2746
rect 2325 2694 2377 2746
rect 2389 2694 2441 2746
rect 2453 2694 2505 2746
rect 2517 2694 2569 2746
rect 4883 2694 4935 2746
rect 4947 2694 4999 2746
rect 5011 2694 5063 2746
rect 5075 2694 5127 2746
rect 5139 2694 5191 2746
rect 7505 2694 7557 2746
rect 7569 2694 7621 2746
rect 7633 2694 7685 2746
rect 7697 2694 7749 2746
rect 7761 2694 7813 2746
rect 10127 2694 10179 2746
rect 10191 2694 10243 2746
rect 10255 2694 10307 2746
rect 10319 2694 10371 2746
rect 10383 2694 10435 2746
rect 2921 2150 2973 2202
rect 2985 2150 3037 2202
rect 3049 2150 3101 2202
rect 3113 2150 3165 2202
rect 3177 2150 3229 2202
rect 5543 2150 5595 2202
rect 5607 2150 5659 2202
rect 5671 2150 5723 2202
rect 5735 2150 5787 2202
rect 5799 2150 5851 2202
rect 8165 2150 8217 2202
rect 8229 2150 8281 2202
rect 8293 2150 8345 2202
rect 8357 2150 8409 2202
rect 8421 2150 8473 2202
rect 10787 2150 10839 2202
rect 10851 2150 10903 2202
rect 10915 2150 10967 2202
rect 10979 2150 11031 2202
rect 11043 2150 11095 2202
<< metal2 >>
rect 2261 12540 2569 12549
rect 2261 12538 2267 12540
rect 2323 12538 2347 12540
rect 2403 12538 2427 12540
rect 2483 12538 2507 12540
rect 2563 12538 2569 12540
rect 2323 12486 2325 12538
rect 2505 12486 2507 12538
rect 2261 12484 2267 12486
rect 2323 12484 2347 12486
rect 2403 12484 2427 12486
rect 2483 12484 2507 12486
rect 2563 12484 2569 12486
rect 2261 12475 2569 12484
rect 4883 12540 5191 12549
rect 4883 12538 4889 12540
rect 4945 12538 4969 12540
rect 5025 12538 5049 12540
rect 5105 12538 5129 12540
rect 5185 12538 5191 12540
rect 4945 12486 4947 12538
rect 5127 12486 5129 12538
rect 4883 12484 4889 12486
rect 4945 12484 4969 12486
rect 5025 12484 5049 12486
rect 5105 12484 5129 12486
rect 5185 12484 5191 12486
rect 4883 12475 5191 12484
rect 7505 12540 7813 12549
rect 7505 12538 7511 12540
rect 7567 12538 7591 12540
rect 7647 12538 7671 12540
rect 7727 12538 7751 12540
rect 7807 12538 7813 12540
rect 7567 12486 7569 12538
rect 7749 12486 7751 12538
rect 7505 12484 7511 12486
rect 7567 12484 7591 12486
rect 7647 12484 7671 12486
rect 7727 12484 7751 12486
rect 7807 12484 7813 12486
rect 7505 12475 7813 12484
rect 10127 12540 10435 12549
rect 10127 12538 10133 12540
rect 10189 12538 10213 12540
rect 10269 12538 10293 12540
rect 10349 12538 10373 12540
rect 10429 12538 10435 12540
rect 10189 12486 10191 12538
rect 10371 12486 10373 12538
rect 10127 12484 10133 12486
rect 10189 12484 10213 12486
rect 10269 12484 10293 12486
rect 10349 12484 10373 12486
rect 10429 12484 10435 12486
rect 10127 12475 10435 12484
rect 2921 11996 3229 12005
rect 2921 11994 2927 11996
rect 2983 11994 3007 11996
rect 3063 11994 3087 11996
rect 3143 11994 3167 11996
rect 3223 11994 3229 11996
rect 2983 11942 2985 11994
rect 3165 11942 3167 11994
rect 2921 11940 2927 11942
rect 2983 11940 3007 11942
rect 3063 11940 3087 11942
rect 3143 11940 3167 11942
rect 3223 11940 3229 11942
rect 2921 11931 3229 11940
rect 5543 11996 5851 12005
rect 5543 11994 5549 11996
rect 5605 11994 5629 11996
rect 5685 11994 5709 11996
rect 5765 11994 5789 11996
rect 5845 11994 5851 11996
rect 5605 11942 5607 11994
rect 5787 11942 5789 11994
rect 5543 11940 5549 11942
rect 5605 11940 5629 11942
rect 5685 11940 5709 11942
rect 5765 11940 5789 11942
rect 5845 11940 5851 11942
rect 5543 11931 5851 11940
rect 8165 11996 8473 12005
rect 8165 11994 8171 11996
rect 8227 11994 8251 11996
rect 8307 11994 8331 11996
rect 8387 11994 8411 11996
rect 8467 11994 8473 11996
rect 8227 11942 8229 11994
rect 8409 11942 8411 11994
rect 8165 11940 8171 11942
rect 8227 11940 8251 11942
rect 8307 11940 8331 11942
rect 8387 11940 8411 11942
rect 8467 11940 8473 11942
rect 8165 11931 8473 11940
rect 10787 11996 11095 12005
rect 10787 11994 10793 11996
rect 10849 11994 10873 11996
rect 10929 11994 10953 11996
rect 11009 11994 11033 11996
rect 11089 11994 11095 11996
rect 10849 11942 10851 11994
rect 11031 11942 11033 11994
rect 10787 11940 10793 11942
rect 10849 11940 10873 11942
rect 10929 11940 10953 11942
rect 11009 11940 11033 11942
rect 11089 11940 11095 11942
rect 10787 11931 11095 11940
rect 2261 11452 2569 11461
rect 2261 11450 2267 11452
rect 2323 11450 2347 11452
rect 2403 11450 2427 11452
rect 2483 11450 2507 11452
rect 2563 11450 2569 11452
rect 2323 11398 2325 11450
rect 2505 11398 2507 11450
rect 2261 11396 2267 11398
rect 2323 11396 2347 11398
rect 2403 11396 2427 11398
rect 2483 11396 2507 11398
rect 2563 11396 2569 11398
rect 2261 11387 2569 11396
rect 4883 11452 5191 11461
rect 4883 11450 4889 11452
rect 4945 11450 4969 11452
rect 5025 11450 5049 11452
rect 5105 11450 5129 11452
rect 5185 11450 5191 11452
rect 4945 11398 4947 11450
rect 5127 11398 5129 11450
rect 4883 11396 4889 11398
rect 4945 11396 4969 11398
rect 5025 11396 5049 11398
rect 5105 11396 5129 11398
rect 5185 11396 5191 11398
rect 4883 11387 5191 11396
rect 7505 11452 7813 11461
rect 7505 11450 7511 11452
rect 7567 11450 7591 11452
rect 7647 11450 7671 11452
rect 7727 11450 7751 11452
rect 7807 11450 7813 11452
rect 7567 11398 7569 11450
rect 7749 11398 7751 11450
rect 7505 11396 7511 11398
rect 7567 11396 7591 11398
rect 7647 11396 7671 11398
rect 7727 11396 7751 11398
rect 7807 11396 7813 11398
rect 7505 11387 7813 11396
rect 10127 11452 10435 11461
rect 10127 11450 10133 11452
rect 10189 11450 10213 11452
rect 10269 11450 10293 11452
rect 10349 11450 10373 11452
rect 10429 11450 10435 11452
rect 10189 11398 10191 11450
rect 10371 11398 10373 11450
rect 10127 11396 10133 11398
rect 10189 11396 10213 11398
rect 10269 11396 10293 11398
rect 10349 11396 10373 11398
rect 10429 11396 10435 11398
rect 10127 11387 10435 11396
rect 2921 10908 3229 10917
rect 2921 10906 2927 10908
rect 2983 10906 3007 10908
rect 3063 10906 3087 10908
rect 3143 10906 3167 10908
rect 3223 10906 3229 10908
rect 2983 10854 2985 10906
rect 3165 10854 3167 10906
rect 2921 10852 2927 10854
rect 2983 10852 3007 10854
rect 3063 10852 3087 10854
rect 3143 10852 3167 10854
rect 3223 10852 3229 10854
rect 2921 10843 3229 10852
rect 5543 10908 5851 10917
rect 5543 10906 5549 10908
rect 5605 10906 5629 10908
rect 5685 10906 5709 10908
rect 5765 10906 5789 10908
rect 5845 10906 5851 10908
rect 5605 10854 5607 10906
rect 5787 10854 5789 10906
rect 5543 10852 5549 10854
rect 5605 10852 5629 10854
rect 5685 10852 5709 10854
rect 5765 10852 5789 10854
rect 5845 10852 5851 10854
rect 5543 10843 5851 10852
rect 8165 10908 8473 10917
rect 8165 10906 8171 10908
rect 8227 10906 8251 10908
rect 8307 10906 8331 10908
rect 8387 10906 8411 10908
rect 8467 10906 8473 10908
rect 8227 10854 8229 10906
rect 8409 10854 8411 10906
rect 8165 10852 8171 10854
rect 8227 10852 8251 10854
rect 8307 10852 8331 10854
rect 8387 10852 8411 10854
rect 8467 10852 8473 10854
rect 8165 10843 8473 10852
rect 10787 10908 11095 10917
rect 10787 10906 10793 10908
rect 10849 10906 10873 10908
rect 10929 10906 10953 10908
rect 11009 10906 11033 10908
rect 11089 10906 11095 10908
rect 10849 10854 10851 10906
rect 11031 10854 11033 10906
rect 10787 10852 10793 10854
rect 10849 10852 10873 10854
rect 10929 10852 10953 10854
rect 11009 10852 11033 10854
rect 11089 10852 11095 10854
rect 10787 10843 11095 10852
rect 2261 10364 2569 10373
rect 2261 10362 2267 10364
rect 2323 10362 2347 10364
rect 2403 10362 2427 10364
rect 2483 10362 2507 10364
rect 2563 10362 2569 10364
rect 2323 10310 2325 10362
rect 2505 10310 2507 10362
rect 2261 10308 2267 10310
rect 2323 10308 2347 10310
rect 2403 10308 2427 10310
rect 2483 10308 2507 10310
rect 2563 10308 2569 10310
rect 2261 10299 2569 10308
rect 4883 10364 5191 10373
rect 4883 10362 4889 10364
rect 4945 10362 4969 10364
rect 5025 10362 5049 10364
rect 5105 10362 5129 10364
rect 5185 10362 5191 10364
rect 4945 10310 4947 10362
rect 5127 10310 5129 10362
rect 4883 10308 4889 10310
rect 4945 10308 4969 10310
rect 5025 10308 5049 10310
rect 5105 10308 5129 10310
rect 5185 10308 5191 10310
rect 4883 10299 5191 10308
rect 7505 10364 7813 10373
rect 7505 10362 7511 10364
rect 7567 10362 7591 10364
rect 7647 10362 7671 10364
rect 7727 10362 7751 10364
rect 7807 10362 7813 10364
rect 7567 10310 7569 10362
rect 7749 10310 7751 10362
rect 7505 10308 7511 10310
rect 7567 10308 7591 10310
rect 7647 10308 7671 10310
rect 7727 10308 7751 10310
rect 7807 10308 7813 10310
rect 7505 10299 7813 10308
rect 10127 10364 10435 10373
rect 10127 10362 10133 10364
rect 10189 10362 10213 10364
rect 10269 10362 10293 10364
rect 10349 10362 10373 10364
rect 10429 10362 10435 10364
rect 10189 10310 10191 10362
rect 10371 10310 10373 10362
rect 10127 10308 10133 10310
rect 10189 10308 10213 10310
rect 10269 10308 10293 10310
rect 10349 10308 10373 10310
rect 10429 10308 10435 10310
rect 10127 10299 10435 10308
rect 2921 9820 3229 9829
rect 2921 9818 2927 9820
rect 2983 9818 3007 9820
rect 3063 9818 3087 9820
rect 3143 9818 3167 9820
rect 3223 9818 3229 9820
rect 2983 9766 2985 9818
rect 3165 9766 3167 9818
rect 2921 9764 2927 9766
rect 2983 9764 3007 9766
rect 3063 9764 3087 9766
rect 3143 9764 3167 9766
rect 3223 9764 3229 9766
rect 2921 9755 3229 9764
rect 5543 9820 5851 9829
rect 5543 9818 5549 9820
rect 5605 9818 5629 9820
rect 5685 9818 5709 9820
rect 5765 9818 5789 9820
rect 5845 9818 5851 9820
rect 5605 9766 5607 9818
rect 5787 9766 5789 9818
rect 5543 9764 5549 9766
rect 5605 9764 5629 9766
rect 5685 9764 5709 9766
rect 5765 9764 5789 9766
rect 5845 9764 5851 9766
rect 5543 9755 5851 9764
rect 8165 9820 8473 9829
rect 8165 9818 8171 9820
rect 8227 9818 8251 9820
rect 8307 9818 8331 9820
rect 8387 9818 8411 9820
rect 8467 9818 8473 9820
rect 8227 9766 8229 9818
rect 8409 9766 8411 9818
rect 8165 9764 8171 9766
rect 8227 9764 8251 9766
rect 8307 9764 8331 9766
rect 8387 9764 8411 9766
rect 8467 9764 8473 9766
rect 8165 9755 8473 9764
rect 10787 9820 11095 9829
rect 10787 9818 10793 9820
rect 10849 9818 10873 9820
rect 10929 9818 10953 9820
rect 11009 9818 11033 9820
rect 11089 9818 11095 9820
rect 10849 9766 10851 9818
rect 11031 9766 11033 9818
rect 10787 9764 10793 9766
rect 10849 9764 10873 9766
rect 10929 9764 10953 9766
rect 11009 9764 11033 9766
rect 11089 9764 11095 9766
rect 10787 9755 11095 9764
rect 2261 9276 2569 9285
rect 2261 9274 2267 9276
rect 2323 9274 2347 9276
rect 2403 9274 2427 9276
rect 2483 9274 2507 9276
rect 2563 9274 2569 9276
rect 2323 9222 2325 9274
rect 2505 9222 2507 9274
rect 2261 9220 2267 9222
rect 2323 9220 2347 9222
rect 2403 9220 2427 9222
rect 2483 9220 2507 9222
rect 2563 9220 2569 9222
rect 2261 9211 2569 9220
rect 4883 9276 5191 9285
rect 4883 9274 4889 9276
rect 4945 9274 4969 9276
rect 5025 9274 5049 9276
rect 5105 9274 5129 9276
rect 5185 9274 5191 9276
rect 4945 9222 4947 9274
rect 5127 9222 5129 9274
rect 4883 9220 4889 9222
rect 4945 9220 4969 9222
rect 5025 9220 5049 9222
rect 5105 9220 5129 9222
rect 5185 9220 5191 9222
rect 4883 9211 5191 9220
rect 7505 9276 7813 9285
rect 7505 9274 7511 9276
rect 7567 9274 7591 9276
rect 7647 9274 7671 9276
rect 7727 9274 7751 9276
rect 7807 9274 7813 9276
rect 7567 9222 7569 9274
rect 7749 9222 7751 9274
rect 7505 9220 7511 9222
rect 7567 9220 7591 9222
rect 7647 9220 7671 9222
rect 7727 9220 7751 9222
rect 7807 9220 7813 9222
rect 7505 9211 7813 9220
rect 10127 9276 10435 9285
rect 10127 9274 10133 9276
rect 10189 9274 10213 9276
rect 10269 9274 10293 9276
rect 10349 9274 10373 9276
rect 10429 9274 10435 9276
rect 10189 9222 10191 9274
rect 10371 9222 10373 9274
rect 10127 9220 10133 9222
rect 10189 9220 10213 9222
rect 10269 9220 10293 9222
rect 10349 9220 10373 9222
rect 10429 9220 10435 9222
rect 10127 9211 10435 9220
rect 2921 8732 3229 8741
rect 2921 8730 2927 8732
rect 2983 8730 3007 8732
rect 3063 8730 3087 8732
rect 3143 8730 3167 8732
rect 3223 8730 3229 8732
rect 2983 8678 2985 8730
rect 3165 8678 3167 8730
rect 2921 8676 2927 8678
rect 2983 8676 3007 8678
rect 3063 8676 3087 8678
rect 3143 8676 3167 8678
rect 3223 8676 3229 8678
rect 2921 8667 3229 8676
rect 5543 8732 5851 8741
rect 5543 8730 5549 8732
rect 5605 8730 5629 8732
rect 5685 8730 5709 8732
rect 5765 8730 5789 8732
rect 5845 8730 5851 8732
rect 5605 8678 5607 8730
rect 5787 8678 5789 8730
rect 5543 8676 5549 8678
rect 5605 8676 5629 8678
rect 5685 8676 5709 8678
rect 5765 8676 5789 8678
rect 5845 8676 5851 8678
rect 5543 8667 5851 8676
rect 8165 8732 8473 8741
rect 8165 8730 8171 8732
rect 8227 8730 8251 8732
rect 8307 8730 8331 8732
rect 8387 8730 8411 8732
rect 8467 8730 8473 8732
rect 8227 8678 8229 8730
rect 8409 8678 8411 8730
rect 8165 8676 8171 8678
rect 8227 8676 8251 8678
rect 8307 8676 8331 8678
rect 8387 8676 8411 8678
rect 8467 8676 8473 8678
rect 8165 8667 8473 8676
rect 10787 8732 11095 8741
rect 10787 8730 10793 8732
rect 10849 8730 10873 8732
rect 10929 8730 10953 8732
rect 11009 8730 11033 8732
rect 11089 8730 11095 8732
rect 10849 8678 10851 8730
rect 11031 8678 11033 8730
rect 10787 8676 10793 8678
rect 10849 8676 10873 8678
rect 10929 8676 10953 8678
rect 11009 8676 11033 8678
rect 11089 8676 11095 8678
rect 10787 8667 11095 8676
rect 2261 8188 2569 8197
rect 2261 8186 2267 8188
rect 2323 8186 2347 8188
rect 2403 8186 2427 8188
rect 2483 8186 2507 8188
rect 2563 8186 2569 8188
rect 2323 8134 2325 8186
rect 2505 8134 2507 8186
rect 2261 8132 2267 8134
rect 2323 8132 2347 8134
rect 2403 8132 2427 8134
rect 2483 8132 2507 8134
rect 2563 8132 2569 8134
rect 2261 8123 2569 8132
rect 4883 8188 5191 8197
rect 4883 8186 4889 8188
rect 4945 8186 4969 8188
rect 5025 8186 5049 8188
rect 5105 8186 5129 8188
rect 5185 8186 5191 8188
rect 4945 8134 4947 8186
rect 5127 8134 5129 8186
rect 4883 8132 4889 8134
rect 4945 8132 4969 8134
rect 5025 8132 5049 8134
rect 5105 8132 5129 8134
rect 5185 8132 5191 8134
rect 4883 8123 5191 8132
rect 7505 8188 7813 8197
rect 7505 8186 7511 8188
rect 7567 8186 7591 8188
rect 7647 8186 7671 8188
rect 7727 8186 7751 8188
rect 7807 8186 7813 8188
rect 7567 8134 7569 8186
rect 7749 8134 7751 8186
rect 7505 8132 7511 8134
rect 7567 8132 7591 8134
rect 7647 8132 7671 8134
rect 7727 8132 7751 8134
rect 7807 8132 7813 8134
rect 7505 8123 7813 8132
rect 10127 8188 10435 8197
rect 10127 8186 10133 8188
rect 10189 8186 10213 8188
rect 10269 8186 10293 8188
rect 10349 8186 10373 8188
rect 10429 8186 10435 8188
rect 10189 8134 10191 8186
rect 10371 8134 10373 8186
rect 10127 8132 10133 8134
rect 10189 8132 10213 8134
rect 10269 8132 10293 8134
rect 10349 8132 10373 8134
rect 10429 8132 10435 8134
rect 10127 8123 10435 8132
rect 848 7880 900 7886
rect 848 7822 900 7828
rect 7196 7880 7248 7886
rect 7196 7822 7248 7828
rect 860 7721 888 7822
rect 1584 7744 1636 7750
rect 846 7712 902 7721
rect 1584 7686 1636 7692
rect 846 7647 902 7656
rect 1596 7410 1624 7686
rect 2921 7644 3229 7653
rect 2921 7642 2927 7644
rect 2983 7642 3007 7644
rect 3063 7642 3087 7644
rect 3143 7642 3167 7644
rect 3223 7642 3229 7644
rect 2983 7590 2985 7642
rect 3165 7590 3167 7642
rect 2921 7588 2927 7590
rect 2983 7588 3007 7590
rect 3063 7588 3087 7590
rect 3143 7588 3167 7590
rect 3223 7588 3229 7590
rect 2921 7579 3229 7588
rect 5543 7644 5851 7653
rect 5543 7642 5549 7644
rect 5605 7642 5629 7644
rect 5685 7642 5709 7644
rect 5765 7642 5789 7644
rect 5845 7642 5851 7644
rect 5605 7590 5607 7642
rect 5787 7590 5789 7642
rect 5543 7588 5549 7590
rect 5605 7588 5629 7590
rect 5685 7588 5709 7590
rect 5765 7588 5789 7590
rect 5845 7588 5851 7590
rect 5543 7579 5851 7588
rect 7208 7546 7236 7822
rect 11244 7744 11296 7750
rect 11244 7686 11296 7692
rect 8165 7644 8473 7653
rect 8165 7642 8171 7644
rect 8227 7642 8251 7644
rect 8307 7642 8331 7644
rect 8387 7642 8411 7644
rect 8467 7642 8473 7644
rect 8227 7590 8229 7642
rect 8409 7590 8411 7642
rect 8165 7588 8171 7590
rect 8227 7588 8251 7590
rect 8307 7588 8331 7590
rect 8387 7588 8411 7590
rect 8467 7588 8473 7590
rect 8165 7579 8473 7588
rect 10787 7644 11095 7653
rect 10787 7642 10793 7644
rect 10849 7642 10873 7644
rect 10929 7642 10953 7644
rect 11009 7642 11033 7644
rect 11089 7642 11095 7644
rect 10849 7590 10851 7642
rect 11031 7590 11033 7642
rect 10787 7588 10793 7590
rect 10849 7588 10873 7590
rect 10929 7588 10953 7590
rect 11009 7588 11033 7590
rect 11089 7588 11095 7590
rect 10787 7579 11095 7588
rect 11256 7585 11284 7686
rect 11242 7576 11298 7585
rect 7196 7540 7248 7546
rect 11242 7511 11298 7520
rect 7196 7482 7248 7488
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 1412 6905 1440 7346
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 2261 7100 2569 7109
rect 2261 7098 2267 7100
rect 2323 7098 2347 7100
rect 2403 7098 2427 7100
rect 2483 7098 2507 7100
rect 2563 7098 2569 7100
rect 2323 7046 2325 7098
rect 2505 7046 2507 7098
rect 2261 7044 2267 7046
rect 2323 7044 2347 7046
rect 2403 7044 2427 7046
rect 2483 7044 2507 7046
rect 2563 7044 2569 7046
rect 2261 7035 2569 7044
rect 4883 7100 5191 7109
rect 4883 7098 4889 7100
rect 4945 7098 4969 7100
rect 5025 7098 5049 7100
rect 5105 7098 5129 7100
rect 5185 7098 5191 7100
rect 4945 7046 4947 7098
rect 5127 7046 5129 7098
rect 4883 7044 4889 7046
rect 4945 7044 4969 7046
rect 5025 7044 5049 7046
rect 5105 7044 5129 7046
rect 5185 7044 5191 7046
rect 4883 7035 5191 7044
rect 7505 7100 7813 7109
rect 7505 7098 7511 7100
rect 7567 7098 7591 7100
rect 7647 7098 7671 7100
rect 7727 7098 7751 7100
rect 7807 7098 7813 7100
rect 7567 7046 7569 7098
rect 7749 7046 7751 7098
rect 7505 7044 7511 7046
rect 7567 7044 7591 7046
rect 7647 7044 7671 7046
rect 7727 7044 7751 7046
rect 7807 7044 7813 7046
rect 7505 7035 7813 7044
rect 10127 7100 10435 7109
rect 10127 7098 10133 7100
rect 10189 7098 10213 7100
rect 10269 7098 10293 7100
rect 10349 7098 10373 7100
rect 10429 7098 10435 7100
rect 10189 7046 10191 7098
rect 10371 7046 10373 7098
rect 10127 7044 10133 7046
rect 10189 7044 10213 7046
rect 10269 7044 10293 7046
rect 10349 7044 10373 7046
rect 10429 7044 10435 7046
rect 10127 7035 10435 7044
rect 11164 6905 11192 7142
rect 1398 6896 1454 6905
rect 1398 6831 1454 6840
rect 11150 6896 11206 6905
rect 11150 6831 11206 6840
rect 2921 6556 3229 6565
rect 2921 6554 2927 6556
rect 2983 6554 3007 6556
rect 3063 6554 3087 6556
rect 3143 6554 3167 6556
rect 3223 6554 3229 6556
rect 2983 6502 2985 6554
rect 3165 6502 3167 6554
rect 2921 6500 2927 6502
rect 2983 6500 3007 6502
rect 3063 6500 3087 6502
rect 3143 6500 3167 6502
rect 3223 6500 3229 6502
rect 2921 6491 3229 6500
rect 5543 6556 5851 6565
rect 5543 6554 5549 6556
rect 5605 6554 5629 6556
rect 5685 6554 5709 6556
rect 5765 6554 5789 6556
rect 5845 6554 5851 6556
rect 5605 6502 5607 6554
rect 5787 6502 5789 6554
rect 5543 6500 5549 6502
rect 5605 6500 5629 6502
rect 5685 6500 5709 6502
rect 5765 6500 5789 6502
rect 5845 6500 5851 6502
rect 5543 6491 5851 6500
rect 8165 6556 8473 6565
rect 8165 6554 8171 6556
rect 8227 6554 8251 6556
rect 8307 6554 8331 6556
rect 8387 6554 8411 6556
rect 8467 6554 8473 6556
rect 8227 6502 8229 6554
rect 8409 6502 8411 6554
rect 8165 6500 8171 6502
rect 8227 6500 8251 6502
rect 8307 6500 8331 6502
rect 8387 6500 8411 6502
rect 8467 6500 8473 6502
rect 8165 6491 8473 6500
rect 10787 6556 11095 6565
rect 10787 6554 10793 6556
rect 10849 6554 10873 6556
rect 10929 6554 10953 6556
rect 11009 6554 11033 6556
rect 11089 6554 11095 6556
rect 10849 6502 10851 6554
rect 11031 6502 11033 6554
rect 10787 6500 10793 6502
rect 10849 6500 10873 6502
rect 10929 6500 10953 6502
rect 11009 6500 11033 6502
rect 11089 6500 11095 6502
rect 10787 6491 11095 6500
rect 2261 6012 2569 6021
rect 2261 6010 2267 6012
rect 2323 6010 2347 6012
rect 2403 6010 2427 6012
rect 2483 6010 2507 6012
rect 2563 6010 2569 6012
rect 2323 5958 2325 6010
rect 2505 5958 2507 6010
rect 2261 5956 2267 5958
rect 2323 5956 2347 5958
rect 2403 5956 2427 5958
rect 2483 5956 2507 5958
rect 2563 5956 2569 5958
rect 2261 5947 2569 5956
rect 4883 6012 5191 6021
rect 4883 6010 4889 6012
rect 4945 6010 4969 6012
rect 5025 6010 5049 6012
rect 5105 6010 5129 6012
rect 5185 6010 5191 6012
rect 4945 5958 4947 6010
rect 5127 5958 5129 6010
rect 4883 5956 4889 5958
rect 4945 5956 4969 5958
rect 5025 5956 5049 5958
rect 5105 5956 5129 5958
rect 5185 5956 5191 5958
rect 4883 5947 5191 5956
rect 7505 6012 7813 6021
rect 7505 6010 7511 6012
rect 7567 6010 7591 6012
rect 7647 6010 7671 6012
rect 7727 6010 7751 6012
rect 7807 6010 7813 6012
rect 7567 5958 7569 6010
rect 7749 5958 7751 6010
rect 7505 5956 7511 5958
rect 7567 5956 7591 5958
rect 7647 5956 7671 5958
rect 7727 5956 7751 5958
rect 7807 5956 7813 5958
rect 7505 5947 7813 5956
rect 10127 6012 10435 6021
rect 10127 6010 10133 6012
rect 10189 6010 10213 6012
rect 10269 6010 10293 6012
rect 10349 6010 10373 6012
rect 10429 6010 10435 6012
rect 10189 5958 10191 6010
rect 10371 5958 10373 6010
rect 10127 5956 10133 5958
rect 10189 5956 10213 5958
rect 10269 5956 10293 5958
rect 10349 5956 10373 5958
rect 10429 5956 10435 5958
rect 10127 5947 10435 5956
rect 2921 5468 3229 5477
rect 2921 5466 2927 5468
rect 2983 5466 3007 5468
rect 3063 5466 3087 5468
rect 3143 5466 3167 5468
rect 3223 5466 3229 5468
rect 2983 5414 2985 5466
rect 3165 5414 3167 5466
rect 2921 5412 2927 5414
rect 2983 5412 3007 5414
rect 3063 5412 3087 5414
rect 3143 5412 3167 5414
rect 3223 5412 3229 5414
rect 2921 5403 3229 5412
rect 5543 5468 5851 5477
rect 5543 5466 5549 5468
rect 5605 5466 5629 5468
rect 5685 5466 5709 5468
rect 5765 5466 5789 5468
rect 5845 5466 5851 5468
rect 5605 5414 5607 5466
rect 5787 5414 5789 5466
rect 5543 5412 5549 5414
rect 5605 5412 5629 5414
rect 5685 5412 5709 5414
rect 5765 5412 5789 5414
rect 5845 5412 5851 5414
rect 5543 5403 5851 5412
rect 8165 5468 8473 5477
rect 8165 5466 8171 5468
rect 8227 5466 8251 5468
rect 8307 5466 8331 5468
rect 8387 5466 8411 5468
rect 8467 5466 8473 5468
rect 8227 5414 8229 5466
rect 8409 5414 8411 5466
rect 8165 5412 8171 5414
rect 8227 5412 8251 5414
rect 8307 5412 8331 5414
rect 8387 5412 8411 5414
rect 8467 5412 8473 5414
rect 8165 5403 8473 5412
rect 10787 5468 11095 5477
rect 10787 5466 10793 5468
rect 10849 5466 10873 5468
rect 10929 5466 10953 5468
rect 11009 5466 11033 5468
rect 11089 5466 11095 5468
rect 10849 5414 10851 5466
rect 11031 5414 11033 5466
rect 10787 5412 10793 5414
rect 10849 5412 10873 5414
rect 10929 5412 10953 5414
rect 11009 5412 11033 5414
rect 11089 5412 11095 5414
rect 10787 5403 11095 5412
rect 2261 4924 2569 4933
rect 2261 4922 2267 4924
rect 2323 4922 2347 4924
rect 2403 4922 2427 4924
rect 2483 4922 2507 4924
rect 2563 4922 2569 4924
rect 2323 4870 2325 4922
rect 2505 4870 2507 4922
rect 2261 4868 2267 4870
rect 2323 4868 2347 4870
rect 2403 4868 2427 4870
rect 2483 4868 2507 4870
rect 2563 4868 2569 4870
rect 2261 4859 2569 4868
rect 4883 4924 5191 4933
rect 4883 4922 4889 4924
rect 4945 4922 4969 4924
rect 5025 4922 5049 4924
rect 5105 4922 5129 4924
rect 5185 4922 5191 4924
rect 4945 4870 4947 4922
rect 5127 4870 5129 4922
rect 4883 4868 4889 4870
rect 4945 4868 4969 4870
rect 5025 4868 5049 4870
rect 5105 4868 5129 4870
rect 5185 4868 5191 4870
rect 4883 4859 5191 4868
rect 7505 4924 7813 4933
rect 7505 4922 7511 4924
rect 7567 4922 7591 4924
rect 7647 4922 7671 4924
rect 7727 4922 7751 4924
rect 7807 4922 7813 4924
rect 7567 4870 7569 4922
rect 7749 4870 7751 4922
rect 7505 4868 7511 4870
rect 7567 4868 7591 4870
rect 7647 4868 7671 4870
rect 7727 4868 7751 4870
rect 7807 4868 7813 4870
rect 7505 4859 7813 4868
rect 10127 4924 10435 4933
rect 10127 4922 10133 4924
rect 10189 4922 10213 4924
rect 10269 4922 10293 4924
rect 10349 4922 10373 4924
rect 10429 4922 10435 4924
rect 10189 4870 10191 4922
rect 10371 4870 10373 4922
rect 10127 4868 10133 4870
rect 10189 4868 10213 4870
rect 10269 4868 10293 4870
rect 10349 4868 10373 4870
rect 10429 4868 10435 4870
rect 10127 4859 10435 4868
rect 2921 4380 3229 4389
rect 2921 4378 2927 4380
rect 2983 4378 3007 4380
rect 3063 4378 3087 4380
rect 3143 4378 3167 4380
rect 3223 4378 3229 4380
rect 2983 4326 2985 4378
rect 3165 4326 3167 4378
rect 2921 4324 2927 4326
rect 2983 4324 3007 4326
rect 3063 4324 3087 4326
rect 3143 4324 3167 4326
rect 3223 4324 3229 4326
rect 2921 4315 3229 4324
rect 5543 4380 5851 4389
rect 5543 4378 5549 4380
rect 5605 4378 5629 4380
rect 5685 4378 5709 4380
rect 5765 4378 5789 4380
rect 5845 4378 5851 4380
rect 5605 4326 5607 4378
rect 5787 4326 5789 4378
rect 5543 4324 5549 4326
rect 5605 4324 5629 4326
rect 5685 4324 5709 4326
rect 5765 4324 5789 4326
rect 5845 4324 5851 4326
rect 5543 4315 5851 4324
rect 8165 4380 8473 4389
rect 8165 4378 8171 4380
rect 8227 4378 8251 4380
rect 8307 4378 8331 4380
rect 8387 4378 8411 4380
rect 8467 4378 8473 4380
rect 8227 4326 8229 4378
rect 8409 4326 8411 4378
rect 8165 4324 8171 4326
rect 8227 4324 8251 4326
rect 8307 4324 8331 4326
rect 8387 4324 8411 4326
rect 8467 4324 8473 4326
rect 8165 4315 8473 4324
rect 10787 4380 11095 4389
rect 10787 4378 10793 4380
rect 10849 4378 10873 4380
rect 10929 4378 10953 4380
rect 11009 4378 11033 4380
rect 11089 4378 11095 4380
rect 10849 4326 10851 4378
rect 11031 4326 11033 4378
rect 10787 4324 10793 4326
rect 10849 4324 10873 4326
rect 10929 4324 10953 4326
rect 11009 4324 11033 4326
rect 11089 4324 11095 4326
rect 10787 4315 11095 4324
rect 2261 3836 2569 3845
rect 2261 3834 2267 3836
rect 2323 3834 2347 3836
rect 2403 3834 2427 3836
rect 2483 3834 2507 3836
rect 2563 3834 2569 3836
rect 2323 3782 2325 3834
rect 2505 3782 2507 3834
rect 2261 3780 2267 3782
rect 2323 3780 2347 3782
rect 2403 3780 2427 3782
rect 2483 3780 2507 3782
rect 2563 3780 2569 3782
rect 2261 3771 2569 3780
rect 4883 3836 5191 3845
rect 4883 3834 4889 3836
rect 4945 3834 4969 3836
rect 5025 3834 5049 3836
rect 5105 3834 5129 3836
rect 5185 3834 5191 3836
rect 4945 3782 4947 3834
rect 5127 3782 5129 3834
rect 4883 3780 4889 3782
rect 4945 3780 4969 3782
rect 5025 3780 5049 3782
rect 5105 3780 5129 3782
rect 5185 3780 5191 3782
rect 4883 3771 5191 3780
rect 7505 3836 7813 3845
rect 7505 3834 7511 3836
rect 7567 3834 7591 3836
rect 7647 3834 7671 3836
rect 7727 3834 7751 3836
rect 7807 3834 7813 3836
rect 7567 3782 7569 3834
rect 7749 3782 7751 3834
rect 7505 3780 7511 3782
rect 7567 3780 7591 3782
rect 7647 3780 7671 3782
rect 7727 3780 7751 3782
rect 7807 3780 7813 3782
rect 7505 3771 7813 3780
rect 10127 3836 10435 3845
rect 10127 3834 10133 3836
rect 10189 3834 10213 3836
rect 10269 3834 10293 3836
rect 10349 3834 10373 3836
rect 10429 3834 10435 3836
rect 10189 3782 10191 3834
rect 10371 3782 10373 3834
rect 10127 3780 10133 3782
rect 10189 3780 10213 3782
rect 10269 3780 10293 3782
rect 10349 3780 10373 3782
rect 10429 3780 10435 3782
rect 10127 3771 10435 3780
rect 2921 3292 3229 3301
rect 2921 3290 2927 3292
rect 2983 3290 3007 3292
rect 3063 3290 3087 3292
rect 3143 3290 3167 3292
rect 3223 3290 3229 3292
rect 2983 3238 2985 3290
rect 3165 3238 3167 3290
rect 2921 3236 2927 3238
rect 2983 3236 3007 3238
rect 3063 3236 3087 3238
rect 3143 3236 3167 3238
rect 3223 3236 3229 3238
rect 2921 3227 3229 3236
rect 5543 3292 5851 3301
rect 5543 3290 5549 3292
rect 5605 3290 5629 3292
rect 5685 3290 5709 3292
rect 5765 3290 5789 3292
rect 5845 3290 5851 3292
rect 5605 3238 5607 3290
rect 5787 3238 5789 3290
rect 5543 3236 5549 3238
rect 5605 3236 5629 3238
rect 5685 3236 5709 3238
rect 5765 3236 5789 3238
rect 5845 3236 5851 3238
rect 5543 3227 5851 3236
rect 8165 3292 8473 3301
rect 8165 3290 8171 3292
rect 8227 3290 8251 3292
rect 8307 3290 8331 3292
rect 8387 3290 8411 3292
rect 8467 3290 8473 3292
rect 8227 3238 8229 3290
rect 8409 3238 8411 3290
rect 8165 3236 8171 3238
rect 8227 3236 8251 3238
rect 8307 3236 8331 3238
rect 8387 3236 8411 3238
rect 8467 3236 8473 3238
rect 8165 3227 8473 3236
rect 10787 3292 11095 3301
rect 10787 3290 10793 3292
rect 10849 3290 10873 3292
rect 10929 3290 10953 3292
rect 11009 3290 11033 3292
rect 11089 3290 11095 3292
rect 10849 3238 10851 3290
rect 11031 3238 11033 3290
rect 10787 3236 10793 3238
rect 10849 3236 10873 3238
rect 10929 3236 10953 3238
rect 11009 3236 11033 3238
rect 11089 3236 11095 3238
rect 10787 3227 11095 3236
rect 2261 2748 2569 2757
rect 2261 2746 2267 2748
rect 2323 2746 2347 2748
rect 2403 2746 2427 2748
rect 2483 2746 2507 2748
rect 2563 2746 2569 2748
rect 2323 2694 2325 2746
rect 2505 2694 2507 2746
rect 2261 2692 2267 2694
rect 2323 2692 2347 2694
rect 2403 2692 2427 2694
rect 2483 2692 2507 2694
rect 2563 2692 2569 2694
rect 2261 2683 2569 2692
rect 4883 2748 5191 2757
rect 4883 2746 4889 2748
rect 4945 2746 4969 2748
rect 5025 2746 5049 2748
rect 5105 2746 5129 2748
rect 5185 2746 5191 2748
rect 4945 2694 4947 2746
rect 5127 2694 5129 2746
rect 4883 2692 4889 2694
rect 4945 2692 4969 2694
rect 5025 2692 5049 2694
rect 5105 2692 5129 2694
rect 5185 2692 5191 2694
rect 4883 2683 5191 2692
rect 7505 2748 7813 2757
rect 7505 2746 7511 2748
rect 7567 2746 7591 2748
rect 7647 2746 7671 2748
rect 7727 2746 7751 2748
rect 7807 2746 7813 2748
rect 7567 2694 7569 2746
rect 7749 2694 7751 2746
rect 7505 2692 7511 2694
rect 7567 2692 7591 2694
rect 7647 2692 7671 2694
rect 7727 2692 7751 2694
rect 7807 2692 7813 2694
rect 7505 2683 7813 2692
rect 10127 2748 10435 2757
rect 10127 2746 10133 2748
rect 10189 2746 10213 2748
rect 10269 2746 10293 2748
rect 10349 2746 10373 2748
rect 10429 2746 10435 2748
rect 10189 2694 10191 2746
rect 10371 2694 10373 2746
rect 10127 2692 10133 2694
rect 10189 2692 10213 2694
rect 10269 2692 10293 2694
rect 10349 2692 10373 2694
rect 10429 2692 10435 2694
rect 10127 2683 10435 2692
rect 2921 2204 3229 2213
rect 2921 2202 2927 2204
rect 2983 2202 3007 2204
rect 3063 2202 3087 2204
rect 3143 2202 3167 2204
rect 3223 2202 3229 2204
rect 2983 2150 2985 2202
rect 3165 2150 3167 2202
rect 2921 2148 2927 2150
rect 2983 2148 3007 2150
rect 3063 2148 3087 2150
rect 3143 2148 3167 2150
rect 3223 2148 3229 2150
rect 2921 2139 3229 2148
rect 5543 2204 5851 2213
rect 5543 2202 5549 2204
rect 5605 2202 5629 2204
rect 5685 2202 5709 2204
rect 5765 2202 5789 2204
rect 5845 2202 5851 2204
rect 5605 2150 5607 2202
rect 5787 2150 5789 2202
rect 5543 2148 5549 2150
rect 5605 2148 5629 2150
rect 5685 2148 5709 2150
rect 5765 2148 5789 2150
rect 5845 2148 5851 2150
rect 5543 2139 5851 2148
rect 8165 2204 8473 2213
rect 8165 2202 8171 2204
rect 8227 2202 8251 2204
rect 8307 2202 8331 2204
rect 8387 2202 8411 2204
rect 8467 2202 8473 2204
rect 8227 2150 8229 2202
rect 8409 2150 8411 2202
rect 8165 2148 8171 2150
rect 8227 2148 8251 2150
rect 8307 2148 8331 2150
rect 8387 2148 8411 2150
rect 8467 2148 8473 2150
rect 8165 2139 8473 2148
rect 10787 2204 11095 2213
rect 10787 2202 10793 2204
rect 10849 2202 10873 2204
rect 10929 2202 10953 2204
rect 11009 2202 11033 2204
rect 11089 2202 11095 2204
rect 10849 2150 10851 2202
rect 11031 2150 11033 2202
rect 10787 2148 10793 2150
rect 10849 2148 10873 2150
rect 10929 2148 10953 2150
rect 11009 2148 11033 2150
rect 11089 2148 11095 2150
rect 10787 2139 11095 2148
<< via2 >>
rect 2267 12538 2323 12540
rect 2347 12538 2403 12540
rect 2427 12538 2483 12540
rect 2507 12538 2563 12540
rect 2267 12486 2313 12538
rect 2313 12486 2323 12538
rect 2347 12486 2377 12538
rect 2377 12486 2389 12538
rect 2389 12486 2403 12538
rect 2427 12486 2441 12538
rect 2441 12486 2453 12538
rect 2453 12486 2483 12538
rect 2507 12486 2517 12538
rect 2517 12486 2563 12538
rect 2267 12484 2323 12486
rect 2347 12484 2403 12486
rect 2427 12484 2483 12486
rect 2507 12484 2563 12486
rect 4889 12538 4945 12540
rect 4969 12538 5025 12540
rect 5049 12538 5105 12540
rect 5129 12538 5185 12540
rect 4889 12486 4935 12538
rect 4935 12486 4945 12538
rect 4969 12486 4999 12538
rect 4999 12486 5011 12538
rect 5011 12486 5025 12538
rect 5049 12486 5063 12538
rect 5063 12486 5075 12538
rect 5075 12486 5105 12538
rect 5129 12486 5139 12538
rect 5139 12486 5185 12538
rect 4889 12484 4945 12486
rect 4969 12484 5025 12486
rect 5049 12484 5105 12486
rect 5129 12484 5185 12486
rect 7511 12538 7567 12540
rect 7591 12538 7647 12540
rect 7671 12538 7727 12540
rect 7751 12538 7807 12540
rect 7511 12486 7557 12538
rect 7557 12486 7567 12538
rect 7591 12486 7621 12538
rect 7621 12486 7633 12538
rect 7633 12486 7647 12538
rect 7671 12486 7685 12538
rect 7685 12486 7697 12538
rect 7697 12486 7727 12538
rect 7751 12486 7761 12538
rect 7761 12486 7807 12538
rect 7511 12484 7567 12486
rect 7591 12484 7647 12486
rect 7671 12484 7727 12486
rect 7751 12484 7807 12486
rect 10133 12538 10189 12540
rect 10213 12538 10269 12540
rect 10293 12538 10349 12540
rect 10373 12538 10429 12540
rect 10133 12486 10179 12538
rect 10179 12486 10189 12538
rect 10213 12486 10243 12538
rect 10243 12486 10255 12538
rect 10255 12486 10269 12538
rect 10293 12486 10307 12538
rect 10307 12486 10319 12538
rect 10319 12486 10349 12538
rect 10373 12486 10383 12538
rect 10383 12486 10429 12538
rect 10133 12484 10189 12486
rect 10213 12484 10269 12486
rect 10293 12484 10349 12486
rect 10373 12484 10429 12486
rect 2927 11994 2983 11996
rect 3007 11994 3063 11996
rect 3087 11994 3143 11996
rect 3167 11994 3223 11996
rect 2927 11942 2973 11994
rect 2973 11942 2983 11994
rect 3007 11942 3037 11994
rect 3037 11942 3049 11994
rect 3049 11942 3063 11994
rect 3087 11942 3101 11994
rect 3101 11942 3113 11994
rect 3113 11942 3143 11994
rect 3167 11942 3177 11994
rect 3177 11942 3223 11994
rect 2927 11940 2983 11942
rect 3007 11940 3063 11942
rect 3087 11940 3143 11942
rect 3167 11940 3223 11942
rect 5549 11994 5605 11996
rect 5629 11994 5685 11996
rect 5709 11994 5765 11996
rect 5789 11994 5845 11996
rect 5549 11942 5595 11994
rect 5595 11942 5605 11994
rect 5629 11942 5659 11994
rect 5659 11942 5671 11994
rect 5671 11942 5685 11994
rect 5709 11942 5723 11994
rect 5723 11942 5735 11994
rect 5735 11942 5765 11994
rect 5789 11942 5799 11994
rect 5799 11942 5845 11994
rect 5549 11940 5605 11942
rect 5629 11940 5685 11942
rect 5709 11940 5765 11942
rect 5789 11940 5845 11942
rect 8171 11994 8227 11996
rect 8251 11994 8307 11996
rect 8331 11994 8387 11996
rect 8411 11994 8467 11996
rect 8171 11942 8217 11994
rect 8217 11942 8227 11994
rect 8251 11942 8281 11994
rect 8281 11942 8293 11994
rect 8293 11942 8307 11994
rect 8331 11942 8345 11994
rect 8345 11942 8357 11994
rect 8357 11942 8387 11994
rect 8411 11942 8421 11994
rect 8421 11942 8467 11994
rect 8171 11940 8227 11942
rect 8251 11940 8307 11942
rect 8331 11940 8387 11942
rect 8411 11940 8467 11942
rect 10793 11994 10849 11996
rect 10873 11994 10929 11996
rect 10953 11994 11009 11996
rect 11033 11994 11089 11996
rect 10793 11942 10839 11994
rect 10839 11942 10849 11994
rect 10873 11942 10903 11994
rect 10903 11942 10915 11994
rect 10915 11942 10929 11994
rect 10953 11942 10967 11994
rect 10967 11942 10979 11994
rect 10979 11942 11009 11994
rect 11033 11942 11043 11994
rect 11043 11942 11089 11994
rect 10793 11940 10849 11942
rect 10873 11940 10929 11942
rect 10953 11940 11009 11942
rect 11033 11940 11089 11942
rect 2267 11450 2323 11452
rect 2347 11450 2403 11452
rect 2427 11450 2483 11452
rect 2507 11450 2563 11452
rect 2267 11398 2313 11450
rect 2313 11398 2323 11450
rect 2347 11398 2377 11450
rect 2377 11398 2389 11450
rect 2389 11398 2403 11450
rect 2427 11398 2441 11450
rect 2441 11398 2453 11450
rect 2453 11398 2483 11450
rect 2507 11398 2517 11450
rect 2517 11398 2563 11450
rect 2267 11396 2323 11398
rect 2347 11396 2403 11398
rect 2427 11396 2483 11398
rect 2507 11396 2563 11398
rect 4889 11450 4945 11452
rect 4969 11450 5025 11452
rect 5049 11450 5105 11452
rect 5129 11450 5185 11452
rect 4889 11398 4935 11450
rect 4935 11398 4945 11450
rect 4969 11398 4999 11450
rect 4999 11398 5011 11450
rect 5011 11398 5025 11450
rect 5049 11398 5063 11450
rect 5063 11398 5075 11450
rect 5075 11398 5105 11450
rect 5129 11398 5139 11450
rect 5139 11398 5185 11450
rect 4889 11396 4945 11398
rect 4969 11396 5025 11398
rect 5049 11396 5105 11398
rect 5129 11396 5185 11398
rect 7511 11450 7567 11452
rect 7591 11450 7647 11452
rect 7671 11450 7727 11452
rect 7751 11450 7807 11452
rect 7511 11398 7557 11450
rect 7557 11398 7567 11450
rect 7591 11398 7621 11450
rect 7621 11398 7633 11450
rect 7633 11398 7647 11450
rect 7671 11398 7685 11450
rect 7685 11398 7697 11450
rect 7697 11398 7727 11450
rect 7751 11398 7761 11450
rect 7761 11398 7807 11450
rect 7511 11396 7567 11398
rect 7591 11396 7647 11398
rect 7671 11396 7727 11398
rect 7751 11396 7807 11398
rect 10133 11450 10189 11452
rect 10213 11450 10269 11452
rect 10293 11450 10349 11452
rect 10373 11450 10429 11452
rect 10133 11398 10179 11450
rect 10179 11398 10189 11450
rect 10213 11398 10243 11450
rect 10243 11398 10255 11450
rect 10255 11398 10269 11450
rect 10293 11398 10307 11450
rect 10307 11398 10319 11450
rect 10319 11398 10349 11450
rect 10373 11398 10383 11450
rect 10383 11398 10429 11450
rect 10133 11396 10189 11398
rect 10213 11396 10269 11398
rect 10293 11396 10349 11398
rect 10373 11396 10429 11398
rect 2927 10906 2983 10908
rect 3007 10906 3063 10908
rect 3087 10906 3143 10908
rect 3167 10906 3223 10908
rect 2927 10854 2973 10906
rect 2973 10854 2983 10906
rect 3007 10854 3037 10906
rect 3037 10854 3049 10906
rect 3049 10854 3063 10906
rect 3087 10854 3101 10906
rect 3101 10854 3113 10906
rect 3113 10854 3143 10906
rect 3167 10854 3177 10906
rect 3177 10854 3223 10906
rect 2927 10852 2983 10854
rect 3007 10852 3063 10854
rect 3087 10852 3143 10854
rect 3167 10852 3223 10854
rect 5549 10906 5605 10908
rect 5629 10906 5685 10908
rect 5709 10906 5765 10908
rect 5789 10906 5845 10908
rect 5549 10854 5595 10906
rect 5595 10854 5605 10906
rect 5629 10854 5659 10906
rect 5659 10854 5671 10906
rect 5671 10854 5685 10906
rect 5709 10854 5723 10906
rect 5723 10854 5735 10906
rect 5735 10854 5765 10906
rect 5789 10854 5799 10906
rect 5799 10854 5845 10906
rect 5549 10852 5605 10854
rect 5629 10852 5685 10854
rect 5709 10852 5765 10854
rect 5789 10852 5845 10854
rect 8171 10906 8227 10908
rect 8251 10906 8307 10908
rect 8331 10906 8387 10908
rect 8411 10906 8467 10908
rect 8171 10854 8217 10906
rect 8217 10854 8227 10906
rect 8251 10854 8281 10906
rect 8281 10854 8293 10906
rect 8293 10854 8307 10906
rect 8331 10854 8345 10906
rect 8345 10854 8357 10906
rect 8357 10854 8387 10906
rect 8411 10854 8421 10906
rect 8421 10854 8467 10906
rect 8171 10852 8227 10854
rect 8251 10852 8307 10854
rect 8331 10852 8387 10854
rect 8411 10852 8467 10854
rect 10793 10906 10849 10908
rect 10873 10906 10929 10908
rect 10953 10906 11009 10908
rect 11033 10906 11089 10908
rect 10793 10854 10839 10906
rect 10839 10854 10849 10906
rect 10873 10854 10903 10906
rect 10903 10854 10915 10906
rect 10915 10854 10929 10906
rect 10953 10854 10967 10906
rect 10967 10854 10979 10906
rect 10979 10854 11009 10906
rect 11033 10854 11043 10906
rect 11043 10854 11089 10906
rect 10793 10852 10849 10854
rect 10873 10852 10929 10854
rect 10953 10852 11009 10854
rect 11033 10852 11089 10854
rect 2267 10362 2323 10364
rect 2347 10362 2403 10364
rect 2427 10362 2483 10364
rect 2507 10362 2563 10364
rect 2267 10310 2313 10362
rect 2313 10310 2323 10362
rect 2347 10310 2377 10362
rect 2377 10310 2389 10362
rect 2389 10310 2403 10362
rect 2427 10310 2441 10362
rect 2441 10310 2453 10362
rect 2453 10310 2483 10362
rect 2507 10310 2517 10362
rect 2517 10310 2563 10362
rect 2267 10308 2323 10310
rect 2347 10308 2403 10310
rect 2427 10308 2483 10310
rect 2507 10308 2563 10310
rect 4889 10362 4945 10364
rect 4969 10362 5025 10364
rect 5049 10362 5105 10364
rect 5129 10362 5185 10364
rect 4889 10310 4935 10362
rect 4935 10310 4945 10362
rect 4969 10310 4999 10362
rect 4999 10310 5011 10362
rect 5011 10310 5025 10362
rect 5049 10310 5063 10362
rect 5063 10310 5075 10362
rect 5075 10310 5105 10362
rect 5129 10310 5139 10362
rect 5139 10310 5185 10362
rect 4889 10308 4945 10310
rect 4969 10308 5025 10310
rect 5049 10308 5105 10310
rect 5129 10308 5185 10310
rect 7511 10362 7567 10364
rect 7591 10362 7647 10364
rect 7671 10362 7727 10364
rect 7751 10362 7807 10364
rect 7511 10310 7557 10362
rect 7557 10310 7567 10362
rect 7591 10310 7621 10362
rect 7621 10310 7633 10362
rect 7633 10310 7647 10362
rect 7671 10310 7685 10362
rect 7685 10310 7697 10362
rect 7697 10310 7727 10362
rect 7751 10310 7761 10362
rect 7761 10310 7807 10362
rect 7511 10308 7567 10310
rect 7591 10308 7647 10310
rect 7671 10308 7727 10310
rect 7751 10308 7807 10310
rect 10133 10362 10189 10364
rect 10213 10362 10269 10364
rect 10293 10362 10349 10364
rect 10373 10362 10429 10364
rect 10133 10310 10179 10362
rect 10179 10310 10189 10362
rect 10213 10310 10243 10362
rect 10243 10310 10255 10362
rect 10255 10310 10269 10362
rect 10293 10310 10307 10362
rect 10307 10310 10319 10362
rect 10319 10310 10349 10362
rect 10373 10310 10383 10362
rect 10383 10310 10429 10362
rect 10133 10308 10189 10310
rect 10213 10308 10269 10310
rect 10293 10308 10349 10310
rect 10373 10308 10429 10310
rect 2927 9818 2983 9820
rect 3007 9818 3063 9820
rect 3087 9818 3143 9820
rect 3167 9818 3223 9820
rect 2927 9766 2973 9818
rect 2973 9766 2983 9818
rect 3007 9766 3037 9818
rect 3037 9766 3049 9818
rect 3049 9766 3063 9818
rect 3087 9766 3101 9818
rect 3101 9766 3113 9818
rect 3113 9766 3143 9818
rect 3167 9766 3177 9818
rect 3177 9766 3223 9818
rect 2927 9764 2983 9766
rect 3007 9764 3063 9766
rect 3087 9764 3143 9766
rect 3167 9764 3223 9766
rect 5549 9818 5605 9820
rect 5629 9818 5685 9820
rect 5709 9818 5765 9820
rect 5789 9818 5845 9820
rect 5549 9766 5595 9818
rect 5595 9766 5605 9818
rect 5629 9766 5659 9818
rect 5659 9766 5671 9818
rect 5671 9766 5685 9818
rect 5709 9766 5723 9818
rect 5723 9766 5735 9818
rect 5735 9766 5765 9818
rect 5789 9766 5799 9818
rect 5799 9766 5845 9818
rect 5549 9764 5605 9766
rect 5629 9764 5685 9766
rect 5709 9764 5765 9766
rect 5789 9764 5845 9766
rect 8171 9818 8227 9820
rect 8251 9818 8307 9820
rect 8331 9818 8387 9820
rect 8411 9818 8467 9820
rect 8171 9766 8217 9818
rect 8217 9766 8227 9818
rect 8251 9766 8281 9818
rect 8281 9766 8293 9818
rect 8293 9766 8307 9818
rect 8331 9766 8345 9818
rect 8345 9766 8357 9818
rect 8357 9766 8387 9818
rect 8411 9766 8421 9818
rect 8421 9766 8467 9818
rect 8171 9764 8227 9766
rect 8251 9764 8307 9766
rect 8331 9764 8387 9766
rect 8411 9764 8467 9766
rect 10793 9818 10849 9820
rect 10873 9818 10929 9820
rect 10953 9818 11009 9820
rect 11033 9818 11089 9820
rect 10793 9766 10839 9818
rect 10839 9766 10849 9818
rect 10873 9766 10903 9818
rect 10903 9766 10915 9818
rect 10915 9766 10929 9818
rect 10953 9766 10967 9818
rect 10967 9766 10979 9818
rect 10979 9766 11009 9818
rect 11033 9766 11043 9818
rect 11043 9766 11089 9818
rect 10793 9764 10849 9766
rect 10873 9764 10929 9766
rect 10953 9764 11009 9766
rect 11033 9764 11089 9766
rect 2267 9274 2323 9276
rect 2347 9274 2403 9276
rect 2427 9274 2483 9276
rect 2507 9274 2563 9276
rect 2267 9222 2313 9274
rect 2313 9222 2323 9274
rect 2347 9222 2377 9274
rect 2377 9222 2389 9274
rect 2389 9222 2403 9274
rect 2427 9222 2441 9274
rect 2441 9222 2453 9274
rect 2453 9222 2483 9274
rect 2507 9222 2517 9274
rect 2517 9222 2563 9274
rect 2267 9220 2323 9222
rect 2347 9220 2403 9222
rect 2427 9220 2483 9222
rect 2507 9220 2563 9222
rect 4889 9274 4945 9276
rect 4969 9274 5025 9276
rect 5049 9274 5105 9276
rect 5129 9274 5185 9276
rect 4889 9222 4935 9274
rect 4935 9222 4945 9274
rect 4969 9222 4999 9274
rect 4999 9222 5011 9274
rect 5011 9222 5025 9274
rect 5049 9222 5063 9274
rect 5063 9222 5075 9274
rect 5075 9222 5105 9274
rect 5129 9222 5139 9274
rect 5139 9222 5185 9274
rect 4889 9220 4945 9222
rect 4969 9220 5025 9222
rect 5049 9220 5105 9222
rect 5129 9220 5185 9222
rect 7511 9274 7567 9276
rect 7591 9274 7647 9276
rect 7671 9274 7727 9276
rect 7751 9274 7807 9276
rect 7511 9222 7557 9274
rect 7557 9222 7567 9274
rect 7591 9222 7621 9274
rect 7621 9222 7633 9274
rect 7633 9222 7647 9274
rect 7671 9222 7685 9274
rect 7685 9222 7697 9274
rect 7697 9222 7727 9274
rect 7751 9222 7761 9274
rect 7761 9222 7807 9274
rect 7511 9220 7567 9222
rect 7591 9220 7647 9222
rect 7671 9220 7727 9222
rect 7751 9220 7807 9222
rect 10133 9274 10189 9276
rect 10213 9274 10269 9276
rect 10293 9274 10349 9276
rect 10373 9274 10429 9276
rect 10133 9222 10179 9274
rect 10179 9222 10189 9274
rect 10213 9222 10243 9274
rect 10243 9222 10255 9274
rect 10255 9222 10269 9274
rect 10293 9222 10307 9274
rect 10307 9222 10319 9274
rect 10319 9222 10349 9274
rect 10373 9222 10383 9274
rect 10383 9222 10429 9274
rect 10133 9220 10189 9222
rect 10213 9220 10269 9222
rect 10293 9220 10349 9222
rect 10373 9220 10429 9222
rect 2927 8730 2983 8732
rect 3007 8730 3063 8732
rect 3087 8730 3143 8732
rect 3167 8730 3223 8732
rect 2927 8678 2973 8730
rect 2973 8678 2983 8730
rect 3007 8678 3037 8730
rect 3037 8678 3049 8730
rect 3049 8678 3063 8730
rect 3087 8678 3101 8730
rect 3101 8678 3113 8730
rect 3113 8678 3143 8730
rect 3167 8678 3177 8730
rect 3177 8678 3223 8730
rect 2927 8676 2983 8678
rect 3007 8676 3063 8678
rect 3087 8676 3143 8678
rect 3167 8676 3223 8678
rect 5549 8730 5605 8732
rect 5629 8730 5685 8732
rect 5709 8730 5765 8732
rect 5789 8730 5845 8732
rect 5549 8678 5595 8730
rect 5595 8678 5605 8730
rect 5629 8678 5659 8730
rect 5659 8678 5671 8730
rect 5671 8678 5685 8730
rect 5709 8678 5723 8730
rect 5723 8678 5735 8730
rect 5735 8678 5765 8730
rect 5789 8678 5799 8730
rect 5799 8678 5845 8730
rect 5549 8676 5605 8678
rect 5629 8676 5685 8678
rect 5709 8676 5765 8678
rect 5789 8676 5845 8678
rect 8171 8730 8227 8732
rect 8251 8730 8307 8732
rect 8331 8730 8387 8732
rect 8411 8730 8467 8732
rect 8171 8678 8217 8730
rect 8217 8678 8227 8730
rect 8251 8678 8281 8730
rect 8281 8678 8293 8730
rect 8293 8678 8307 8730
rect 8331 8678 8345 8730
rect 8345 8678 8357 8730
rect 8357 8678 8387 8730
rect 8411 8678 8421 8730
rect 8421 8678 8467 8730
rect 8171 8676 8227 8678
rect 8251 8676 8307 8678
rect 8331 8676 8387 8678
rect 8411 8676 8467 8678
rect 10793 8730 10849 8732
rect 10873 8730 10929 8732
rect 10953 8730 11009 8732
rect 11033 8730 11089 8732
rect 10793 8678 10839 8730
rect 10839 8678 10849 8730
rect 10873 8678 10903 8730
rect 10903 8678 10915 8730
rect 10915 8678 10929 8730
rect 10953 8678 10967 8730
rect 10967 8678 10979 8730
rect 10979 8678 11009 8730
rect 11033 8678 11043 8730
rect 11043 8678 11089 8730
rect 10793 8676 10849 8678
rect 10873 8676 10929 8678
rect 10953 8676 11009 8678
rect 11033 8676 11089 8678
rect 2267 8186 2323 8188
rect 2347 8186 2403 8188
rect 2427 8186 2483 8188
rect 2507 8186 2563 8188
rect 2267 8134 2313 8186
rect 2313 8134 2323 8186
rect 2347 8134 2377 8186
rect 2377 8134 2389 8186
rect 2389 8134 2403 8186
rect 2427 8134 2441 8186
rect 2441 8134 2453 8186
rect 2453 8134 2483 8186
rect 2507 8134 2517 8186
rect 2517 8134 2563 8186
rect 2267 8132 2323 8134
rect 2347 8132 2403 8134
rect 2427 8132 2483 8134
rect 2507 8132 2563 8134
rect 4889 8186 4945 8188
rect 4969 8186 5025 8188
rect 5049 8186 5105 8188
rect 5129 8186 5185 8188
rect 4889 8134 4935 8186
rect 4935 8134 4945 8186
rect 4969 8134 4999 8186
rect 4999 8134 5011 8186
rect 5011 8134 5025 8186
rect 5049 8134 5063 8186
rect 5063 8134 5075 8186
rect 5075 8134 5105 8186
rect 5129 8134 5139 8186
rect 5139 8134 5185 8186
rect 4889 8132 4945 8134
rect 4969 8132 5025 8134
rect 5049 8132 5105 8134
rect 5129 8132 5185 8134
rect 7511 8186 7567 8188
rect 7591 8186 7647 8188
rect 7671 8186 7727 8188
rect 7751 8186 7807 8188
rect 7511 8134 7557 8186
rect 7557 8134 7567 8186
rect 7591 8134 7621 8186
rect 7621 8134 7633 8186
rect 7633 8134 7647 8186
rect 7671 8134 7685 8186
rect 7685 8134 7697 8186
rect 7697 8134 7727 8186
rect 7751 8134 7761 8186
rect 7761 8134 7807 8186
rect 7511 8132 7567 8134
rect 7591 8132 7647 8134
rect 7671 8132 7727 8134
rect 7751 8132 7807 8134
rect 10133 8186 10189 8188
rect 10213 8186 10269 8188
rect 10293 8186 10349 8188
rect 10373 8186 10429 8188
rect 10133 8134 10179 8186
rect 10179 8134 10189 8186
rect 10213 8134 10243 8186
rect 10243 8134 10255 8186
rect 10255 8134 10269 8186
rect 10293 8134 10307 8186
rect 10307 8134 10319 8186
rect 10319 8134 10349 8186
rect 10373 8134 10383 8186
rect 10383 8134 10429 8186
rect 10133 8132 10189 8134
rect 10213 8132 10269 8134
rect 10293 8132 10349 8134
rect 10373 8132 10429 8134
rect 846 7656 902 7712
rect 2927 7642 2983 7644
rect 3007 7642 3063 7644
rect 3087 7642 3143 7644
rect 3167 7642 3223 7644
rect 2927 7590 2973 7642
rect 2973 7590 2983 7642
rect 3007 7590 3037 7642
rect 3037 7590 3049 7642
rect 3049 7590 3063 7642
rect 3087 7590 3101 7642
rect 3101 7590 3113 7642
rect 3113 7590 3143 7642
rect 3167 7590 3177 7642
rect 3177 7590 3223 7642
rect 2927 7588 2983 7590
rect 3007 7588 3063 7590
rect 3087 7588 3143 7590
rect 3167 7588 3223 7590
rect 5549 7642 5605 7644
rect 5629 7642 5685 7644
rect 5709 7642 5765 7644
rect 5789 7642 5845 7644
rect 5549 7590 5595 7642
rect 5595 7590 5605 7642
rect 5629 7590 5659 7642
rect 5659 7590 5671 7642
rect 5671 7590 5685 7642
rect 5709 7590 5723 7642
rect 5723 7590 5735 7642
rect 5735 7590 5765 7642
rect 5789 7590 5799 7642
rect 5799 7590 5845 7642
rect 5549 7588 5605 7590
rect 5629 7588 5685 7590
rect 5709 7588 5765 7590
rect 5789 7588 5845 7590
rect 8171 7642 8227 7644
rect 8251 7642 8307 7644
rect 8331 7642 8387 7644
rect 8411 7642 8467 7644
rect 8171 7590 8217 7642
rect 8217 7590 8227 7642
rect 8251 7590 8281 7642
rect 8281 7590 8293 7642
rect 8293 7590 8307 7642
rect 8331 7590 8345 7642
rect 8345 7590 8357 7642
rect 8357 7590 8387 7642
rect 8411 7590 8421 7642
rect 8421 7590 8467 7642
rect 8171 7588 8227 7590
rect 8251 7588 8307 7590
rect 8331 7588 8387 7590
rect 8411 7588 8467 7590
rect 10793 7642 10849 7644
rect 10873 7642 10929 7644
rect 10953 7642 11009 7644
rect 11033 7642 11089 7644
rect 10793 7590 10839 7642
rect 10839 7590 10849 7642
rect 10873 7590 10903 7642
rect 10903 7590 10915 7642
rect 10915 7590 10929 7642
rect 10953 7590 10967 7642
rect 10967 7590 10979 7642
rect 10979 7590 11009 7642
rect 11033 7590 11043 7642
rect 11043 7590 11089 7642
rect 10793 7588 10849 7590
rect 10873 7588 10929 7590
rect 10953 7588 11009 7590
rect 11033 7588 11089 7590
rect 11242 7520 11298 7576
rect 2267 7098 2323 7100
rect 2347 7098 2403 7100
rect 2427 7098 2483 7100
rect 2507 7098 2563 7100
rect 2267 7046 2313 7098
rect 2313 7046 2323 7098
rect 2347 7046 2377 7098
rect 2377 7046 2389 7098
rect 2389 7046 2403 7098
rect 2427 7046 2441 7098
rect 2441 7046 2453 7098
rect 2453 7046 2483 7098
rect 2507 7046 2517 7098
rect 2517 7046 2563 7098
rect 2267 7044 2323 7046
rect 2347 7044 2403 7046
rect 2427 7044 2483 7046
rect 2507 7044 2563 7046
rect 4889 7098 4945 7100
rect 4969 7098 5025 7100
rect 5049 7098 5105 7100
rect 5129 7098 5185 7100
rect 4889 7046 4935 7098
rect 4935 7046 4945 7098
rect 4969 7046 4999 7098
rect 4999 7046 5011 7098
rect 5011 7046 5025 7098
rect 5049 7046 5063 7098
rect 5063 7046 5075 7098
rect 5075 7046 5105 7098
rect 5129 7046 5139 7098
rect 5139 7046 5185 7098
rect 4889 7044 4945 7046
rect 4969 7044 5025 7046
rect 5049 7044 5105 7046
rect 5129 7044 5185 7046
rect 7511 7098 7567 7100
rect 7591 7098 7647 7100
rect 7671 7098 7727 7100
rect 7751 7098 7807 7100
rect 7511 7046 7557 7098
rect 7557 7046 7567 7098
rect 7591 7046 7621 7098
rect 7621 7046 7633 7098
rect 7633 7046 7647 7098
rect 7671 7046 7685 7098
rect 7685 7046 7697 7098
rect 7697 7046 7727 7098
rect 7751 7046 7761 7098
rect 7761 7046 7807 7098
rect 7511 7044 7567 7046
rect 7591 7044 7647 7046
rect 7671 7044 7727 7046
rect 7751 7044 7807 7046
rect 10133 7098 10189 7100
rect 10213 7098 10269 7100
rect 10293 7098 10349 7100
rect 10373 7098 10429 7100
rect 10133 7046 10179 7098
rect 10179 7046 10189 7098
rect 10213 7046 10243 7098
rect 10243 7046 10255 7098
rect 10255 7046 10269 7098
rect 10293 7046 10307 7098
rect 10307 7046 10319 7098
rect 10319 7046 10349 7098
rect 10373 7046 10383 7098
rect 10383 7046 10429 7098
rect 10133 7044 10189 7046
rect 10213 7044 10269 7046
rect 10293 7044 10349 7046
rect 10373 7044 10429 7046
rect 1398 6840 1454 6896
rect 11150 6840 11206 6896
rect 2927 6554 2983 6556
rect 3007 6554 3063 6556
rect 3087 6554 3143 6556
rect 3167 6554 3223 6556
rect 2927 6502 2973 6554
rect 2973 6502 2983 6554
rect 3007 6502 3037 6554
rect 3037 6502 3049 6554
rect 3049 6502 3063 6554
rect 3087 6502 3101 6554
rect 3101 6502 3113 6554
rect 3113 6502 3143 6554
rect 3167 6502 3177 6554
rect 3177 6502 3223 6554
rect 2927 6500 2983 6502
rect 3007 6500 3063 6502
rect 3087 6500 3143 6502
rect 3167 6500 3223 6502
rect 5549 6554 5605 6556
rect 5629 6554 5685 6556
rect 5709 6554 5765 6556
rect 5789 6554 5845 6556
rect 5549 6502 5595 6554
rect 5595 6502 5605 6554
rect 5629 6502 5659 6554
rect 5659 6502 5671 6554
rect 5671 6502 5685 6554
rect 5709 6502 5723 6554
rect 5723 6502 5735 6554
rect 5735 6502 5765 6554
rect 5789 6502 5799 6554
rect 5799 6502 5845 6554
rect 5549 6500 5605 6502
rect 5629 6500 5685 6502
rect 5709 6500 5765 6502
rect 5789 6500 5845 6502
rect 8171 6554 8227 6556
rect 8251 6554 8307 6556
rect 8331 6554 8387 6556
rect 8411 6554 8467 6556
rect 8171 6502 8217 6554
rect 8217 6502 8227 6554
rect 8251 6502 8281 6554
rect 8281 6502 8293 6554
rect 8293 6502 8307 6554
rect 8331 6502 8345 6554
rect 8345 6502 8357 6554
rect 8357 6502 8387 6554
rect 8411 6502 8421 6554
rect 8421 6502 8467 6554
rect 8171 6500 8227 6502
rect 8251 6500 8307 6502
rect 8331 6500 8387 6502
rect 8411 6500 8467 6502
rect 10793 6554 10849 6556
rect 10873 6554 10929 6556
rect 10953 6554 11009 6556
rect 11033 6554 11089 6556
rect 10793 6502 10839 6554
rect 10839 6502 10849 6554
rect 10873 6502 10903 6554
rect 10903 6502 10915 6554
rect 10915 6502 10929 6554
rect 10953 6502 10967 6554
rect 10967 6502 10979 6554
rect 10979 6502 11009 6554
rect 11033 6502 11043 6554
rect 11043 6502 11089 6554
rect 10793 6500 10849 6502
rect 10873 6500 10929 6502
rect 10953 6500 11009 6502
rect 11033 6500 11089 6502
rect 2267 6010 2323 6012
rect 2347 6010 2403 6012
rect 2427 6010 2483 6012
rect 2507 6010 2563 6012
rect 2267 5958 2313 6010
rect 2313 5958 2323 6010
rect 2347 5958 2377 6010
rect 2377 5958 2389 6010
rect 2389 5958 2403 6010
rect 2427 5958 2441 6010
rect 2441 5958 2453 6010
rect 2453 5958 2483 6010
rect 2507 5958 2517 6010
rect 2517 5958 2563 6010
rect 2267 5956 2323 5958
rect 2347 5956 2403 5958
rect 2427 5956 2483 5958
rect 2507 5956 2563 5958
rect 4889 6010 4945 6012
rect 4969 6010 5025 6012
rect 5049 6010 5105 6012
rect 5129 6010 5185 6012
rect 4889 5958 4935 6010
rect 4935 5958 4945 6010
rect 4969 5958 4999 6010
rect 4999 5958 5011 6010
rect 5011 5958 5025 6010
rect 5049 5958 5063 6010
rect 5063 5958 5075 6010
rect 5075 5958 5105 6010
rect 5129 5958 5139 6010
rect 5139 5958 5185 6010
rect 4889 5956 4945 5958
rect 4969 5956 5025 5958
rect 5049 5956 5105 5958
rect 5129 5956 5185 5958
rect 7511 6010 7567 6012
rect 7591 6010 7647 6012
rect 7671 6010 7727 6012
rect 7751 6010 7807 6012
rect 7511 5958 7557 6010
rect 7557 5958 7567 6010
rect 7591 5958 7621 6010
rect 7621 5958 7633 6010
rect 7633 5958 7647 6010
rect 7671 5958 7685 6010
rect 7685 5958 7697 6010
rect 7697 5958 7727 6010
rect 7751 5958 7761 6010
rect 7761 5958 7807 6010
rect 7511 5956 7567 5958
rect 7591 5956 7647 5958
rect 7671 5956 7727 5958
rect 7751 5956 7807 5958
rect 10133 6010 10189 6012
rect 10213 6010 10269 6012
rect 10293 6010 10349 6012
rect 10373 6010 10429 6012
rect 10133 5958 10179 6010
rect 10179 5958 10189 6010
rect 10213 5958 10243 6010
rect 10243 5958 10255 6010
rect 10255 5958 10269 6010
rect 10293 5958 10307 6010
rect 10307 5958 10319 6010
rect 10319 5958 10349 6010
rect 10373 5958 10383 6010
rect 10383 5958 10429 6010
rect 10133 5956 10189 5958
rect 10213 5956 10269 5958
rect 10293 5956 10349 5958
rect 10373 5956 10429 5958
rect 2927 5466 2983 5468
rect 3007 5466 3063 5468
rect 3087 5466 3143 5468
rect 3167 5466 3223 5468
rect 2927 5414 2973 5466
rect 2973 5414 2983 5466
rect 3007 5414 3037 5466
rect 3037 5414 3049 5466
rect 3049 5414 3063 5466
rect 3087 5414 3101 5466
rect 3101 5414 3113 5466
rect 3113 5414 3143 5466
rect 3167 5414 3177 5466
rect 3177 5414 3223 5466
rect 2927 5412 2983 5414
rect 3007 5412 3063 5414
rect 3087 5412 3143 5414
rect 3167 5412 3223 5414
rect 5549 5466 5605 5468
rect 5629 5466 5685 5468
rect 5709 5466 5765 5468
rect 5789 5466 5845 5468
rect 5549 5414 5595 5466
rect 5595 5414 5605 5466
rect 5629 5414 5659 5466
rect 5659 5414 5671 5466
rect 5671 5414 5685 5466
rect 5709 5414 5723 5466
rect 5723 5414 5735 5466
rect 5735 5414 5765 5466
rect 5789 5414 5799 5466
rect 5799 5414 5845 5466
rect 5549 5412 5605 5414
rect 5629 5412 5685 5414
rect 5709 5412 5765 5414
rect 5789 5412 5845 5414
rect 8171 5466 8227 5468
rect 8251 5466 8307 5468
rect 8331 5466 8387 5468
rect 8411 5466 8467 5468
rect 8171 5414 8217 5466
rect 8217 5414 8227 5466
rect 8251 5414 8281 5466
rect 8281 5414 8293 5466
rect 8293 5414 8307 5466
rect 8331 5414 8345 5466
rect 8345 5414 8357 5466
rect 8357 5414 8387 5466
rect 8411 5414 8421 5466
rect 8421 5414 8467 5466
rect 8171 5412 8227 5414
rect 8251 5412 8307 5414
rect 8331 5412 8387 5414
rect 8411 5412 8467 5414
rect 10793 5466 10849 5468
rect 10873 5466 10929 5468
rect 10953 5466 11009 5468
rect 11033 5466 11089 5468
rect 10793 5414 10839 5466
rect 10839 5414 10849 5466
rect 10873 5414 10903 5466
rect 10903 5414 10915 5466
rect 10915 5414 10929 5466
rect 10953 5414 10967 5466
rect 10967 5414 10979 5466
rect 10979 5414 11009 5466
rect 11033 5414 11043 5466
rect 11043 5414 11089 5466
rect 10793 5412 10849 5414
rect 10873 5412 10929 5414
rect 10953 5412 11009 5414
rect 11033 5412 11089 5414
rect 2267 4922 2323 4924
rect 2347 4922 2403 4924
rect 2427 4922 2483 4924
rect 2507 4922 2563 4924
rect 2267 4870 2313 4922
rect 2313 4870 2323 4922
rect 2347 4870 2377 4922
rect 2377 4870 2389 4922
rect 2389 4870 2403 4922
rect 2427 4870 2441 4922
rect 2441 4870 2453 4922
rect 2453 4870 2483 4922
rect 2507 4870 2517 4922
rect 2517 4870 2563 4922
rect 2267 4868 2323 4870
rect 2347 4868 2403 4870
rect 2427 4868 2483 4870
rect 2507 4868 2563 4870
rect 4889 4922 4945 4924
rect 4969 4922 5025 4924
rect 5049 4922 5105 4924
rect 5129 4922 5185 4924
rect 4889 4870 4935 4922
rect 4935 4870 4945 4922
rect 4969 4870 4999 4922
rect 4999 4870 5011 4922
rect 5011 4870 5025 4922
rect 5049 4870 5063 4922
rect 5063 4870 5075 4922
rect 5075 4870 5105 4922
rect 5129 4870 5139 4922
rect 5139 4870 5185 4922
rect 4889 4868 4945 4870
rect 4969 4868 5025 4870
rect 5049 4868 5105 4870
rect 5129 4868 5185 4870
rect 7511 4922 7567 4924
rect 7591 4922 7647 4924
rect 7671 4922 7727 4924
rect 7751 4922 7807 4924
rect 7511 4870 7557 4922
rect 7557 4870 7567 4922
rect 7591 4870 7621 4922
rect 7621 4870 7633 4922
rect 7633 4870 7647 4922
rect 7671 4870 7685 4922
rect 7685 4870 7697 4922
rect 7697 4870 7727 4922
rect 7751 4870 7761 4922
rect 7761 4870 7807 4922
rect 7511 4868 7567 4870
rect 7591 4868 7647 4870
rect 7671 4868 7727 4870
rect 7751 4868 7807 4870
rect 10133 4922 10189 4924
rect 10213 4922 10269 4924
rect 10293 4922 10349 4924
rect 10373 4922 10429 4924
rect 10133 4870 10179 4922
rect 10179 4870 10189 4922
rect 10213 4870 10243 4922
rect 10243 4870 10255 4922
rect 10255 4870 10269 4922
rect 10293 4870 10307 4922
rect 10307 4870 10319 4922
rect 10319 4870 10349 4922
rect 10373 4870 10383 4922
rect 10383 4870 10429 4922
rect 10133 4868 10189 4870
rect 10213 4868 10269 4870
rect 10293 4868 10349 4870
rect 10373 4868 10429 4870
rect 2927 4378 2983 4380
rect 3007 4378 3063 4380
rect 3087 4378 3143 4380
rect 3167 4378 3223 4380
rect 2927 4326 2973 4378
rect 2973 4326 2983 4378
rect 3007 4326 3037 4378
rect 3037 4326 3049 4378
rect 3049 4326 3063 4378
rect 3087 4326 3101 4378
rect 3101 4326 3113 4378
rect 3113 4326 3143 4378
rect 3167 4326 3177 4378
rect 3177 4326 3223 4378
rect 2927 4324 2983 4326
rect 3007 4324 3063 4326
rect 3087 4324 3143 4326
rect 3167 4324 3223 4326
rect 5549 4378 5605 4380
rect 5629 4378 5685 4380
rect 5709 4378 5765 4380
rect 5789 4378 5845 4380
rect 5549 4326 5595 4378
rect 5595 4326 5605 4378
rect 5629 4326 5659 4378
rect 5659 4326 5671 4378
rect 5671 4326 5685 4378
rect 5709 4326 5723 4378
rect 5723 4326 5735 4378
rect 5735 4326 5765 4378
rect 5789 4326 5799 4378
rect 5799 4326 5845 4378
rect 5549 4324 5605 4326
rect 5629 4324 5685 4326
rect 5709 4324 5765 4326
rect 5789 4324 5845 4326
rect 8171 4378 8227 4380
rect 8251 4378 8307 4380
rect 8331 4378 8387 4380
rect 8411 4378 8467 4380
rect 8171 4326 8217 4378
rect 8217 4326 8227 4378
rect 8251 4326 8281 4378
rect 8281 4326 8293 4378
rect 8293 4326 8307 4378
rect 8331 4326 8345 4378
rect 8345 4326 8357 4378
rect 8357 4326 8387 4378
rect 8411 4326 8421 4378
rect 8421 4326 8467 4378
rect 8171 4324 8227 4326
rect 8251 4324 8307 4326
rect 8331 4324 8387 4326
rect 8411 4324 8467 4326
rect 10793 4378 10849 4380
rect 10873 4378 10929 4380
rect 10953 4378 11009 4380
rect 11033 4378 11089 4380
rect 10793 4326 10839 4378
rect 10839 4326 10849 4378
rect 10873 4326 10903 4378
rect 10903 4326 10915 4378
rect 10915 4326 10929 4378
rect 10953 4326 10967 4378
rect 10967 4326 10979 4378
rect 10979 4326 11009 4378
rect 11033 4326 11043 4378
rect 11043 4326 11089 4378
rect 10793 4324 10849 4326
rect 10873 4324 10929 4326
rect 10953 4324 11009 4326
rect 11033 4324 11089 4326
rect 2267 3834 2323 3836
rect 2347 3834 2403 3836
rect 2427 3834 2483 3836
rect 2507 3834 2563 3836
rect 2267 3782 2313 3834
rect 2313 3782 2323 3834
rect 2347 3782 2377 3834
rect 2377 3782 2389 3834
rect 2389 3782 2403 3834
rect 2427 3782 2441 3834
rect 2441 3782 2453 3834
rect 2453 3782 2483 3834
rect 2507 3782 2517 3834
rect 2517 3782 2563 3834
rect 2267 3780 2323 3782
rect 2347 3780 2403 3782
rect 2427 3780 2483 3782
rect 2507 3780 2563 3782
rect 4889 3834 4945 3836
rect 4969 3834 5025 3836
rect 5049 3834 5105 3836
rect 5129 3834 5185 3836
rect 4889 3782 4935 3834
rect 4935 3782 4945 3834
rect 4969 3782 4999 3834
rect 4999 3782 5011 3834
rect 5011 3782 5025 3834
rect 5049 3782 5063 3834
rect 5063 3782 5075 3834
rect 5075 3782 5105 3834
rect 5129 3782 5139 3834
rect 5139 3782 5185 3834
rect 4889 3780 4945 3782
rect 4969 3780 5025 3782
rect 5049 3780 5105 3782
rect 5129 3780 5185 3782
rect 7511 3834 7567 3836
rect 7591 3834 7647 3836
rect 7671 3834 7727 3836
rect 7751 3834 7807 3836
rect 7511 3782 7557 3834
rect 7557 3782 7567 3834
rect 7591 3782 7621 3834
rect 7621 3782 7633 3834
rect 7633 3782 7647 3834
rect 7671 3782 7685 3834
rect 7685 3782 7697 3834
rect 7697 3782 7727 3834
rect 7751 3782 7761 3834
rect 7761 3782 7807 3834
rect 7511 3780 7567 3782
rect 7591 3780 7647 3782
rect 7671 3780 7727 3782
rect 7751 3780 7807 3782
rect 10133 3834 10189 3836
rect 10213 3834 10269 3836
rect 10293 3834 10349 3836
rect 10373 3834 10429 3836
rect 10133 3782 10179 3834
rect 10179 3782 10189 3834
rect 10213 3782 10243 3834
rect 10243 3782 10255 3834
rect 10255 3782 10269 3834
rect 10293 3782 10307 3834
rect 10307 3782 10319 3834
rect 10319 3782 10349 3834
rect 10373 3782 10383 3834
rect 10383 3782 10429 3834
rect 10133 3780 10189 3782
rect 10213 3780 10269 3782
rect 10293 3780 10349 3782
rect 10373 3780 10429 3782
rect 2927 3290 2983 3292
rect 3007 3290 3063 3292
rect 3087 3290 3143 3292
rect 3167 3290 3223 3292
rect 2927 3238 2973 3290
rect 2973 3238 2983 3290
rect 3007 3238 3037 3290
rect 3037 3238 3049 3290
rect 3049 3238 3063 3290
rect 3087 3238 3101 3290
rect 3101 3238 3113 3290
rect 3113 3238 3143 3290
rect 3167 3238 3177 3290
rect 3177 3238 3223 3290
rect 2927 3236 2983 3238
rect 3007 3236 3063 3238
rect 3087 3236 3143 3238
rect 3167 3236 3223 3238
rect 5549 3290 5605 3292
rect 5629 3290 5685 3292
rect 5709 3290 5765 3292
rect 5789 3290 5845 3292
rect 5549 3238 5595 3290
rect 5595 3238 5605 3290
rect 5629 3238 5659 3290
rect 5659 3238 5671 3290
rect 5671 3238 5685 3290
rect 5709 3238 5723 3290
rect 5723 3238 5735 3290
rect 5735 3238 5765 3290
rect 5789 3238 5799 3290
rect 5799 3238 5845 3290
rect 5549 3236 5605 3238
rect 5629 3236 5685 3238
rect 5709 3236 5765 3238
rect 5789 3236 5845 3238
rect 8171 3290 8227 3292
rect 8251 3290 8307 3292
rect 8331 3290 8387 3292
rect 8411 3290 8467 3292
rect 8171 3238 8217 3290
rect 8217 3238 8227 3290
rect 8251 3238 8281 3290
rect 8281 3238 8293 3290
rect 8293 3238 8307 3290
rect 8331 3238 8345 3290
rect 8345 3238 8357 3290
rect 8357 3238 8387 3290
rect 8411 3238 8421 3290
rect 8421 3238 8467 3290
rect 8171 3236 8227 3238
rect 8251 3236 8307 3238
rect 8331 3236 8387 3238
rect 8411 3236 8467 3238
rect 10793 3290 10849 3292
rect 10873 3290 10929 3292
rect 10953 3290 11009 3292
rect 11033 3290 11089 3292
rect 10793 3238 10839 3290
rect 10839 3238 10849 3290
rect 10873 3238 10903 3290
rect 10903 3238 10915 3290
rect 10915 3238 10929 3290
rect 10953 3238 10967 3290
rect 10967 3238 10979 3290
rect 10979 3238 11009 3290
rect 11033 3238 11043 3290
rect 11043 3238 11089 3290
rect 10793 3236 10849 3238
rect 10873 3236 10929 3238
rect 10953 3236 11009 3238
rect 11033 3236 11089 3238
rect 2267 2746 2323 2748
rect 2347 2746 2403 2748
rect 2427 2746 2483 2748
rect 2507 2746 2563 2748
rect 2267 2694 2313 2746
rect 2313 2694 2323 2746
rect 2347 2694 2377 2746
rect 2377 2694 2389 2746
rect 2389 2694 2403 2746
rect 2427 2694 2441 2746
rect 2441 2694 2453 2746
rect 2453 2694 2483 2746
rect 2507 2694 2517 2746
rect 2517 2694 2563 2746
rect 2267 2692 2323 2694
rect 2347 2692 2403 2694
rect 2427 2692 2483 2694
rect 2507 2692 2563 2694
rect 4889 2746 4945 2748
rect 4969 2746 5025 2748
rect 5049 2746 5105 2748
rect 5129 2746 5185 2748
rect 4889 2694 4935 2746
rect 4935 2694 4945 2746
rect 4969 2694 4999 2746
rect 4999 2694 5011 2746
rect 5011 2694 5025 2746
rect 5049 2694 5063 2746
rect 5063 2694 5075 2746
rect 5075 2694 5105 2746
rect 5129 2694 5139 2746
rect 5139 2694 5185 2746
rect 4889 2692 4945 2694
rect 4969 2692 5025 2694
rect 5049 2692 5105 2694
rect 5129 2692 5185 2694
rect 7511 2746 7567 2748
rect 7591 2746 7647 2748
rect 7671 2746 7727 2748
rect 7751 2746 7807 2748
rect 7511 2694 7557 2746
rect 7557 2694 7567 2746
rect 7591 2694 7621 2746
rect 7621 2694 7633 2746
rect 7633 2694 7647 2746
rect 7671 2694 7685 2746
rect 7685 2694 7697 2746
rect 7697 2694 7727 2746
rect 7751 2694 7761 2746
rect 7761 2694 7807 2746
rect 7511 2692 7567 2694
rect 7591 2692 7647 2694
rect 7671 2692 7727 2694
rect 7751 2692 7807 2694
rect 10133 2746 10189 2748
rect 10213 2746 10269 2748
rect 10293 2746 10349 2748
rect 10373 2746 10429 2748
rect 10133 2694 10179 2746
rect 10179 2694 10189 2746
rect 10213 2694 10243 2746
rect 10243 2694 10255 2746
rect 10255 2694 10269 2746
rect 10293 2694 10307 2746
rect 10307 2694 10319 2746
rect 10319 2694 10349 2746
rect 10373 2694 10383 2746
rect 10383 2694 10429 2746
rect 10133 2692 10189 2694
rect 10213 2692 10269 2694
rect 10293 2692 10349 2694
rect 10373 2692 10429 2694
rect 2927 2202 2983 2204
rect 3007 2202 3063 2204
rect 3087 2202 3143 2204
rect 3167 2202 3223 2204
rect 2927 2150 2973 2202
rect 2973 2150 2983 2202
rect 3007 2150 3037 2202
rect 3037 2150 3049 2202
rect 3049 2150 3063 2202
rect 3087 2150 3101 2202
rect 3101 2150 3113 2202
rect 3113 2150 3143 2202
rect 3167 2150 3177 2202
rect 3177 2150 3223 2202
rect 2927 2148 2983 2150
rect 3007 2148 3063 2150
rect 3087 2148 3143 2150
rect 3167 2148 3223 2150
rect 5549 2202 5605 2204
rect 5629 2202 5685 2204
rect 5709 2202 5765 2204
rect 5789 2202 5845 2204
rect 5549 2150 5595 2202
rect 5595 2150 5605 2202
rect 5629 2150 5659 2202
rect 5659 2150 5671 2202
rect 5671 2150 5685 2202
rect 5709 2150 5723 2202
rect 5723 2150 5735 2202
rect 5735 2150 5765 2202
rect 5789 2150 5799 2202
rect 5799 2150 5845 2202
rect 5549 2148 5605 2150
rect 5629 2148 5685 2150
rect 5709 2148 5765 2150
rect 5789 2148 5845 2150
rect 8171 2202 8227 2204
rect 8251 2202 8307 2204
rect 8331 2202 8387 2204
rect 8411 2202 8467 2204
rect 8171 2150 8217 2202
rect 8217 2150 8227 2202
rect 8251 2150 8281 2202
rect 8281 2150 8293 2202
rect 8293 2150 8307 2202
rect 8331 2150 8345 2202
rect 8345 2150 8357 2202
rect 8357 2150 8387 2202
rect 8411 2150 8421 2202
rect 8421 2150 8467 2202
rect 8171 2148 8227 2150
rect 8251 2148 8307 2150
rect 8331 2148 8387 2150
rect 8411 2148 8467 2150
rect 10793 2202 10849 2204
rect 10873 2202 10929 2204
rect 10953 2202 11009 2204
rect 11033 2202 11089 2204
rect 10793 2150 10839 2202
rect 10839 2150 10849 2202
rect 10873 2150 10903 2202
rect 10903 2150 10915 2202
rect 10915 2150 10929 2202
rect 10953 2150 10967 2202
rect 10967 2150 10979 2202
rect 10979 2150 11009 2202
rect 11033 2150 11043 2202
rect 11043 2150 11089 2202
rect 10793 2148 10849 2150
rect 10873 2148 10929 2150
rect 10953 2148 11009 2150
rect 11033 2148 11089 2150
<< metal3 >>
rect 2257 12544 2573 12545
rect 2257 12480 2263 12544
rect 2327 12480 2343 12544
rect 2407 12480 2423 12544
rect 2487 12480 2503 12544
rect 2567 12480 2573 12544
rect 2257 12479 2573 12480
rect 4879 12544 5195 12545
rect 4879 12480 4885 12544
rect 4949 12480 4965 12544
rect 5029 12480 5045 12544
rect 5109 12480 5125 12544
rect 5189 12480 5195 12544
rect 4879 12479 5195 12480
rect 7501 12544 7817 12545
rect 7501 12480 7507 12544
rect 7571 12480 7587 12544
rect 7651 12480 7667 12544
rect 7731 12480 7747 12544
rect 7811 12480 7817 12544
rect 7501 12479 7817 12480
rect 10123 12544 10439 12545
rect 10123 12480 10129 12544
rect 10193 12480 10209 12544
rect 10273 12480 10289 12544
rect 10353 12480 10369 12544
rect 10433 12480 10439 12544
rect 10123 12479 10439 12480
rect 2917 12000 3233 12001
rect 2917 11936 2923 12000
rect 2987 11936 3003 12000
rect 3067 11936 3083 12000
rect 3147 11936 3163 12000
rect 3227 11936 3233 12000
rect 2917 11935 3233 11936
rect 5539 12000 5855 12001
rect 5539 11936 5545 12000
rect 5609 11936 5625 12000
rect 5689 11936 5705 12000
rect 5769 11936 5785 12000
rect 5849 11936 5855 12000
rect 5539 11935 5855 11936
rect 8161 12000 8477 12001
rect 8161 11936 8167 12000
rect 8231 11936 8247 12000
rect 8311 11936 8327 12000
rect 8391 11936 8407 12000
rect 8471 11936 8477 12000
rect 8161 11935 8477 11936
rect 10783 12000 11099 12001
rect 10783 11936 10789 12000
rect 10853 11936 10869 12000
rect 10933 11936 10949 12000
rect 11013 11936 11029 12000
rect 11093 11936 11099 12000
rect 10783 11935 11099 11936
rect 2257 11456 2573 11457
rect 2257 11392 2263 11456
rect 2327 11392 2343 11456
rect 2407 11392 2423 11456
rect 2487 11392 2503 11456
rect 2567 11392 2573 11456
rect 2257 11391 2573 11392
rect 4879 11456 5195 11457
rect 4879 11392 4885 11456
rect 4949 11392 4965 11456
rect 5029 11392 5045 11456
rect 5109 11392 5125 11456
rect 5189 11392 5195 11456
rect 4879 11391 5195 11392
rect 7501 11456 7817 11457
rect 7501 11392 7507 11456
rect 7571 11392 7587 11456
rect 7651 11392 7667 11456
rect 7731 11392 7747 11456
rect 7811 11392 7817 11456
rect 7501 11391 7817 11392
rect 10123 11456 10439 11457
rect 10123 11392 10129 11456
rect 10193 11392 10209 11456
rect 10273 11392 10289 11456
rect 10353 11392 10369 11456
rect 10433 11392 10439 11456
rect 10123 11391 10439 11392
rect 2917 10912 3233 10913
rect 2917 10848 2923 10912
rect 2987 10848 3003 10912
rect 3067 10848 3083 10912
rect 3147 10848 3163 10912
rect 3227 10848 3233 10912
rect 2917 10847 3233 10848
rect 5539 10912 5855 10913
rect 5539 10848 5545 10912
rect 5609 10848 5625 10912
rect 5689 10848 5705 10912
rect 5769 10848 5785 10912
rect 5849 10848 5855 10912
rect 5539 10847 5855 10848
rect 8161 10912 8477 10913
rect 8161 10848 8167 10912
rect 8231 10848 8247 10912
rect 8311 10848 8327 10912
rect 8391 10848 8407 10912
rect 8471 10848 8477 10912
rect 8161 10847 8477 10848
rect 10783 10912 11099 10913
rect 10783 10848 10789 10912
rect 10853 10848 10869 10912
rect 10933 10848 10949 10912
rect 11013 10848 11029 10912
rect 11093 10848 11099 10912
rect 10783 10847 11099 10848
rect 2257 10368 2573 10369
rect 2257 10304 2263 10368
rect 2327 10304 2343 10368
rect 2407 10304 2423 10368
rect 2487 10304 2503 10368
rect 2567 10304 2573 10368
rect 2257 10303 2573 10304
rect 4879 10368 5195 10369
rect 4879 10304 4885 10368
rect 4949 10304 4965 10368
rect 5029 10304 5045 10368
rect 5109 10304 5125 10368
rect 5189 10304 5195 10368
rect 4879 10303 5195 10304
rect 7501 10368 7817 10369
rect 7501 10304 7507 10368
rect 7571 10304 7587 10368
rect 7651 10304 7667 10368
rect 7731 10304 7747 10368
rect 7811 10304 7817 10368
rect 7501 10303 7817 10304
rect 10123 10368 10439 10369
rect 10123 10304 10129 10368
rect 10193 10304 10209 10368
rect 10273 10304 10289 10368
rect 10353 10304 10369 10368
rect 10433 10304 10439 10368
rect 10123 10303 10439 10304
rect 2917 9824 3233 9825
rect 2917 9760 2923 9824
rect 2987 9760 3003 9824
rect 3067 9760 3083 9824
rect 3147 9760 3163 9824
rect 3227 9760 3233 9824
rect 2917 9759 3233 9760
rect 5539 9824 5855 9825
rect 5539 9760 5545 9824
rect 5609 9760 5625 9824
rect 5689 9760 5705 9824
rect 5769 9760 5785 9824
rect 5849 9760 5855 9824
rect 5539 9759 5855 9760
rect 8161 9824 8477 9825
rect 8161 9760 8167 9824
rect 8231 9760 8247 9824
rect 8311 9760 8327 9824
rect 8391 9760 8407 9824
rect 8471 9760 8477 9824
rect 8161 9759 8477 9760
rect 10783 9824 11099 9825
rect 10783 9760 10789 9824
rect 10853 9760 10869 9824
rect 10933 9760 10949 9824
rect 11013 9760 11029 9824
rect 11093 9760 11099 9824
rect 10783 9759 11099 9760
rect 2257 9280 2573 9281
rect 2257 9216 2263 9280
rect 2327 9216 2343 9280
rect 2407 9216 2423 9280
rect 2487 9216 2503 9280
rect 2567 9216 2573 9280
rect 2257 9215 2573 9216
rect 4879 9280 5195 9281
rect 4879 9216 4885 9280
rect 4949 9216 4965 9280
rect 5029 9216 5045 9280
rect 5109 9216 5125 9280
rect 5189 9216 5195 9280
rect 4879 9215 5195 9216
rect 7501 9280 7817 9281
rect 7501 9216 7507 9280
rect 7571 9216 7587 9280
rect 7651 9216 7667 9280
rect 7731 9216 7747 9280
rect 7811 9216 7817 9280
rect 7501 9215 7817 9216
rect 10123 9280 10439 9281
rect 10123 9216 10129 9280
rect 10193 9216 10209 9280
rect 10273 9216 10289 9280
rect 10353 9216 10369 9280
rect 10433 9216 10439 9280
rect 10123 9215 10439 9216
rect 2917 8736 3233 8737
rect 2917 8672 2923 8736
rect 2987 8672 3003 8736
rect 3067 8672 3083 8736
rect 3147 8672 3163 8736
rect 3227 8672 3233 8736
rect 2917 8671 3233 8672
rect 5539 8736 5855 8737
rect 5539 8672 5545 8736
rect 5609 8672 5625 8736
rect 5689 8672 5705 8736
rect 5769 8672 5785 8736
rect 5849 8672 5855 8736
rect 5539 8671 5855 8672
rect 8161 8736 8477 8737
rect 8161 8672 8167 8736
rect 8231 8672 8247 8736
rect 8311 8672 8327 8736
rect 8391 8672 8407 8736
rect 8471 8672 8477 8736
rect 8161 8671 8477 8672
rect 10783 8736 11099 8737
rect 10783 8672 10789 8736
rect 10853 8672 10869 8736
rect 10933 8672 10949 8736
rect 11013 8672 11029 8736
rect 11093 8672 11099 8736
rect 10783 8671 11099 8672
rect 2257 8192 2573 8193
rect 2257 8128 2263 8192
rect 2327 8128 2343 8192
rect 2407 8128 2423 8192
rect 2487 8128 2503 8192
rect 2567 8128 2573 8192
rect 2257 8127 2573 8128
rect 4879 8192 5195 8193
rect 4879 8128 4885 8192
rect 4949 8128 4965 8192
rect 5029 8128 5045 8192
rect 5109 8128 5125 8192
rect 5189 8128 5195 8192
rect 4879 8127 5195 8128
rect 7501 8192 7817 8193
rect 7501 8128 7507 8192
rect 7571 8128 7587 8192
rect 7651 8128 7667 8192
rect 7731 8128 7747 8192
rect 7811 8128 7817 8192
rect 7501 8127 7817 8128
rect 10123 8192 10439 8193
rect 10123 8128 10129 8192
rect 10193 8128 10209 8192
rect 10273 8128 10289 8192
rect 10353 8128 10369 8192
rect 10433 8128 10439 8192
rect 10123 8127 10439 8128
rect 841 7714 907 7717
rect 798 7712 907 7714
rect 798 7656 846 7712
rect 902 7656 907 7712
rect 798 7651 907 7656
rect 798 7608 858 7651
rect 0 7518 858 7608
rect 2917 7648 3233 7649
rect 2917 7584 2923 7648
rect 2987 7584 3003 7648
rect 3067 7584 3083 7648
rect 3147 7584 3163 7648
rect 3227 7584 3233 7648
rect 2917 7583 3233 7584
rect 5539 7648 5855 7649
rect 5539 7584 5545 7648
rect 5609 7584 5625 7648
rect 5689 7584 5705 7648
rect 5769 7584 5785 7648
rect 5849 7584 5855 7648
rect 5539 7583 5855 7584
rect 8161 7648 8477 7649
rect 8161 7584 8167 7648
rect 8231 7584 8247 7648
rect 8311 7584 8327 7648
rect 8391 7584 8407 7648
rect 8471 7584 8477 7648
rect 8161 7583 8477 7584
rect 10783 7648 11099 7649
rect 10783 7584 10789 7648
rect 10853 7584 10869 7648
rect 10933 7584 10949 7648
rect 11013 7584 11029 7648
rect 11093 7584 11099 7648
rect 10783 7583 11099 7584
rect 11237 7578 11303 7581
rect 11901 7578 12701 7608
rect 11237 7576 12701 7578
rect 11237 7520 11242 7576
rect 11298 7520 12701 7576
rect 11237 7518 12701 7520
rect 0 7488 800 7518
rect 11237 7515 11303 7518
rect 11901 7488 12701 7518
rect 2257 7104 2573 7105
rect 2257 7040 2263 7104
rect 2327 7040 2343 7104
rect 2407 7040 2423 7104
rect 2487 7040 2503 7104
rect 2567 7040 2573 7104
rect 2257 7039 2573 7040
rect 4879 7104 5195 7105
rect 4879 7040 4885 7104
rect 4949 7040 4965 7104
rect 5029 7040 5045 7104
rect 5109 7040 5125 7104
rect 5189 7040 5195 7104
rect 4879 7039 5195 7040
rect 7501 7104 7817 7105
rect 7501 7040 7507 7104
rect 7571 7040 7587 7104
rect 7651 7040 7667 7104
rect 7731 7040 7747 7104
rect 7811 7040 7817 7104
rect 7501 7039 7817 7040
rect 10123 7104 10439 7105
rect 10123 7040 10129 7104
rect 10193 7040 10209 7104
rect 10273 7040 10289 7104
rect 10353 7040 10369 7104
rect 10433 7040 10439 7104
rect 10123 7039 10439 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 11145 6898 11211 6901
rect 11901 6898 12701 6928
rect 11145 6896 12701 6898
rect 11145 6840 11150 6896
rect 11206 6840 12701 6896
rect 11145 6838 12701 6840
rect 11145 6835 11211 6838
rect 11901 6808 12701 6838
rect 2917 6560 3233 6561
rect 2917 6496 2923 6560
rect 2987 6496 3003 6560
rect 3067 6496 3083 6560
rect 3147 6496 3163 6560
rect 3227 6496 3233 6560
rect 2917 6495 3233 6496
rect 5539 6560 5855 6561
rect 5539 6496 5545 6560
rect 5609 6496 5625 6560
rect 5689 6496 5705 6560
rect 5769 6496 5785 6560
rect 5849 6496 5855 6560
rect 5539 6495 5855 6496
rect 8161 6560 8477 6561
rect 8161 6496 8167 6560
rect 8231 6496 8247 6560
rect 8311 6496 8327 6560
rect 8391 6496 8407 6560
rect 8471 6496 8477 6560
rect 8161 6495 8477 6496
rect 10783 6560 11099 6561
rect 10783 6496 10789 6560
rect 10853 6496 10869 6560
rect 10933 6496 10949 6560
rect 11013 6496 11029 6560
rect 11093 6496 11099 6560
rect 10783 6495 11099 6496
rect 2257 6016 2573 6017
rect 2257 5952 2263 6016
rect 2327 5952 2343 6016
rect 2407 5952 2423 6016
rect 2487 5952 2503 6016
rect 2567 5952 2573 6016
rect 2257 5951 2573 5952
rect 4879 6016 5195 6017
rect 4879 5952 4885 6016
rect 4949 5952 4965 6016
rect 5029 5952 5045 6016
rect 5109 5952 5125 6016
rect 5189 5952 5195 6016
rect 4879 5951 5195 5952
rect 7501 6016 7817 6017
rect 7501 5952 7507 6016
rect 7571 5952 7587 6016
rect 7651 5952 7667 6016
rect 7731 5952 7747 6016
rect 7811 5952 7817 6016
rect 7501 5951 7817 5952
rect 10123 6016 10439 6017
rect 10123 5952 10129 6016
rect 10193 5952 10209 6016
rect 10273 5952 10289 6016
rect 10353 5952 10369 6016
rect 10433 5952 10439 6016
rect 10123 5951 10439 5952
rect 2917 5472 3233 5473
rect 2917 5408 2923 5472
rect 2987 5408 3003 5472
rect 3067 5408 3083 5472
rect 3147 5408 3163 5472
rect 3227 5408 3233 5472
rect 2917 5407 3233 5408
rect 5539 5472 5855 5473
rect 5539 5408 5545 5472
rect 5609 5408 5625 5472
rect 5689 5408 5705 5472
rect 5769 5408 5785 5472
rect 5849 5408 5855 5472
rect 5539 5407 5855 5408
rect 8161 5472 8477 5473
rect 8161 5408 8167 5472
rect 8231 5408 8247 5472
rect 8311 5408 8327 5472
rect 8391 5408 8407 5472
rect 8471 5408 8477 5472
rect 8161 5407 8477 5408
rect 10783 5472 11099 5473
rect 10783 5408 10789 5472
rect 10853 5408 10869 5472
rect 10933 5408 10949 5472
rect 11013 5408 11029 5472
rect 11093 5408 11099 5472
rect 10783 5407 11099 5408
rect 2257 4928 2573 4929
rect 2257 4864 2263 4928
rect 2327 4864 2343 4928
rect 2407 4864 2423 4928
rect 2487 4864 2503 4928
rect 2567 4864 2573 4928
rect 2257 4863 2573 4864
rect 4879 4928 5195 4929
rect 4879 4864 4885 4928
rect 4949 4864 4965 4928
rect 5029 4864 5045 4928
rect 5109 4864 5125 4928
rect 5189 4864 5195 4928
rect 4879 4863 5195 4864
rect 7501 4928 7817 4929
rect 7501 4864 7507 4928
rect 7571 4864 7587 4928
rect 7651 4864 7667 4928
rect 7731 4864 7747 4928
rect 7811 4864 7817 4928
rect 7501 4863 7817 4864
rect 10123 4928 10439 4929
rect 10123 4864 10129 4928
rect 10193 4864 10209 4928
rect 10273 4864 10289 4928
rect 10353 4864 10369 4928
rect 10433 4864 10439 4928
rect 10123 4863 10439 4864
rect 2917 4384 3233 4385
rect 2917 4320 2923 4384
rect 2987 4320 3003 4384
rect 3067 4320 3083 4384
rect 3147 4320 3163 4384
rect 3227 4320 3233 4384
rect 2917 4319 3233 4320
rect 5539 4384 5855 4385
rect 5539 4320 5545 4384
rect 5609 4320 5625 4384
rect 5689 4320 5705 4384
rect 5769 4320 5785 4384
rect 5849 4320 5855 4384
rect 5539 4319 5855 4320
rect 8161 4384 8477 4385
rect 8161 4320 8167 4384
rect 8231 4320 8247 4384
rect 8311 4320 8327 4384
rect 8391 4320 8407 4384
rect 8471 4320 8477 4384
rect 8161 4319 8477 4320
rect 10783 4384 11099 4385
rect 10783 4320 10789 4384
rect 10853 4320 10869 4384
rect 10933 4320 10949 4384
rect 11013 4320 11029 4384
rect 11093 4320 11099 4384
rect 10783 4319 11099 4320
rect 2257 3840 2573 3841
rect 2257 3776 2263 3840
rect 2327 3776 2343 3840
rect 2407 3776 2423 3840
rect 2487 3776 2503 3840
rect 2567 3776 2573 3840
rect 2257 3775 2573 3776
rect 4879 3840 5195 3841
rect 4879 3776 4885 3840
rect 4949 3776 4965 3840
rect 5029 3776 5045 3840
rect 5109 3776 5125 3840
rect 5189 3776 5195 3840
rect 4879 3775 5195 3776
rect 7501 3840 7817 3841
rect 7501 3776 7507 3840
rect 7571 3776 7587 3840
rect 7651 3776 7667 3840
rect 7731 3776 7747 3840
rect 7811 3776 7817 3840
rect 7501 3775 7817 3776
rect 10123 3840 10439 3841
rect 10123 3776 10129 3840
rect 10193 3776 10209 3840
rect 10273 3776 10289 3840
rect 10353 3776 10369 3840
rect 10433 3776 10439 3840
rect 10123 3775 10439 3776
rect 2917 3296 3233 3297
rect 2917 3232 2923 3296
rect 2987 3232 3003 3296
rect 3067 3232 3083 3296
rect 3147 3232 3163 3296
rect 3227 3232 3233 3296
rect 2917 3231 3233 3232
rect 5539 3296 5855 3297
rect 5539 3232 5545 3296
rect 5609 3232 5625 3296
rect 5689 3232 5705 3296
rect 5769 3232 5785 3296
rect 5849 3232 5855 3296
rect 5539 3231 5855 3232
rect 8161 3296 8477 3297
rect 8161 3232 8167 3296
rect 8231 3232 8247 3296
rect 8311 3232 8327 3296
rect 8391 3232 8407 3296
rect 8471 3232 8477 3296
rect 8161 3231 8477 3232
rect 10783 3296 11099 3297
rect 10783 3232 10789 3296
rect 10853 3232 10869 3296
rect 10933 3232 10949 3296
rect 11013 3232 11029 3296
rect 11093 3232 11099 3296
rect 10783 3231 11099 3232
rect 2257 2752 2573 2753
rect 2257 2688 2263 2752
rect 2327 2688 2343 2752
rect 2407 2688 2423 2752
rect 2487 2688 2503 2752
rect 2567 2688 2573 2752
rect 2257 2687 2573 2688
rect 4879 2752 5195 2753
rect 4879 2688 4885 2752
rect 4949 2688 4965 2752
rect 5029 2688 5045 2752
rect 5109 2688 5125 2752
rect 5189 2688 5195 2752
rect 4879 2687 5195 2688
rect 7501 2752 7817 2753
rect 7501 2688 7507 2752
rect 7571 2688 7587 2752
rect 7651 2688 7667 2752
rect 7731 2688 7747 2752
rect 7811 2688 7817 2752
rect 7501 2687 7817 2688
rect 10123 2752 10439 2753
rect 10123 2688 10129 2752
rect 10193 2688 10209 2752
rect 10273 2688 10289 2752
rect 10353 2688 10369 2752
rect 10433 2688 10439 2752
rect 10123 2687 10439 2688
rect 2917 2208 3233 2209
rect 2917 2144 2923 2208
rect 2987 2144 3003 2208
rect 3067 2144 3083 2208
rect 3147 2144 3163 2208
rect 3227 2144 3233 2208
rect 2917 2143 3233 2144
rect 5539 2208 5855 2209
rect 5539 2144 5545 2208
rect 5609 2144 5625 2208
rect 5689 2144 5705 2208
rect 5769 2144 5785 2208
rect 5849 2144 5855 2208
rect 5539 2143 5855 2144
rect 8161 2208 8477 2209
rect 8161 2144 8167 2208
rect 8231 2144 8247 2208
rect 8311 2144 8327 2208
rect 8391 2144 8407 2208
rect 8471 2144 8477 2208
rect 8161 2143 8477 2144
rect 10783 2208 11099 2209
rect 10783 2144 10789 2208
rect 10853 2144 10869 2208
rect 10933 2144 10949 2208
rect 11013 2144 11029 2208
rect 11093 2144 11099 2208
rect 10783 2143 11099 2144
<< via3 >>
rect 2263 12540 2327 12544
rect 2263 12484 2267 12540
rect 2267 12484 2323 12540
rect 2323 12484 2327 12540
rect 2263 12480 2327 12484
rect 2343 12540 2407 12544
rect 2343 12484 2347 12540
rect 2347 12484 2403 12540
rect 2403 12484 2407 12540
rect 2343 12480 2407 12484
rect 2423 12540 2487 12544
rect 2423 12484 2427 12540
rect 2427 12484 2483 12540
rect 2483 12484 2487 12540
rect 2423 12480 2487 12484
rect 2503 12540 2567 12544
rect 2503 12484 2507 12540
rect 2507 12484 2563 12540
rect 2563 12484 2567 12540
rect 2503 12480 2567 12484
rect 4885 12540 4949 12544
rect 4885 12484 4889 12540
rect 4889 12484 4945 12540
rect 4945 12484 4949 12540
rect 4885 12480 4949 12484
rect 4965 12540 5029 12544
rect 4965 12484 4969 12540
rect 4969 12484 5025 12540
rect 5025 12484 5029 12540
rect 4965 12480 5029 12484
rect 5045 12540 5109 12544
rect 5045 12484 5049 12540
rect 5049 12484 5105 12540
rect 5105 12484 5109 12540
rect 5045 12480 5109 12484
rect 5125 12540 5189 12544
rect 5125 12484 5129 12540
rect 5129 12484 5185 12540
rect 5185 12484 5189 12540
rect 5125 12480 5189 12484
rect 7507 12540 7571 12544
rect 7507 12484 7511 12540
rect 7511 12484 7567 12540
rect 7567 12484 7571 12540
rect 7507 12480 7571 12484
rect 7587 12540 7651 12544
rect 7587 12484 7591 12540
rect 7591 12484 7647 12540
rect 7647 12484 7651 12540
rect 7587 12480 7651 12484
rect 7667 12540 7731 12544
rect 7667 12484 7671 12540
rect 7671 12484 7727 12540
rect 7727 12484 7731 12540
rect 7667 12480 7731 12484
rect 7747 12540 7811 12544
rect 7747 12484 7751 12540
rect 7751 12484 7807 12540
rect 7807 12484 7811 12540
rect 7747 12480 7811 12484
rect 10129 12540 10193 12544
rect 10129 12484 10133 12540
rect 10133 12484 10189 12540
rect 10189 12484 10193 12540
rect 10129 12480 10193 12484
rect 10209 12540 10273 12544
rect 10209 12484 10213 12540
rect 10213 12484 10269 12540
rect 10269 12484 10273 12540
rect 10209 12480 10273 12484
rect 10289 12540 10353 12544
rect 10289 12484 10293 12540
rect 10293 12484 10349 12540
rect 10349 12484 10353 12540
rect 10289 12480 10353 12484
rect 10369 12540 10433 12544
rect 10369 12484 10373 12540
rect 10373 12484 10429 12540
rect 10429 12484 10433 12540
rect 10369 12480 10433 12484
rect 2923 11996 2987 12000
rect 2923 11940 2927 11996
rect 2927 11940 2983 11996
rect 2983 11940 2987 11996
rect 2923 11936 2987 11940
rect 3003 11996 3067 12000
rect 3003 11940 3007 11996
rect 3007 11940 3063 11996
rect 3063 11940 3067 11996
rect 3003 11936 3067 11940
rect 3083 11996 3147 12000
rect 3083 11940 3087 11996
rect 3087 11940 3143 11996
rect 3143 11940 3147 11996
rect 3083 11936 3147 11940
rect 3163 11996 3227 12000
rect 3163 11940 3167 11996
rect 3167 11940 3223 11996
rect 3223 11940 3227 11996
rect 3163 11936 3227 11940
rect 5545 11996 5609 12000
rect 5545 11940 5549 11996
rect 5549 11940 5605 11996
rect 5605 11940 5609 11996
rect 5545 11936 5609 11940
rect 5625 11996 5689 12000
rect 5625 11940 5629 11996
rect 5629 11940 5685 11996
rect 5685 11940 5689 11996
rect 5625 11936 5689 11940
rect 5705 11996 5769 12000
rect 5705 11940 5709 11996
rect 5709 11940 5765 11996
rect 5765 11940 5769 11996
rect 5705 11936 5769 11940
rect 5785 11996 5849 12000
rect 5785 11940 5789 11996
rect 5789 11940 5845 11996
rect 5845 11940 5849 11996
rect 5785 11936 5849 11940
rect 8167 11996 8231 12000
rect 8167 11940 8171 11996
rect 8171 11940 8227 11996
rect 8227 11940 8231 11996
rect 8167 11936 8231 11940
rect 8247 11996 8311 12000
rect 8247 11940 8251 11996
rect 8251 11940 8307 11996
rect 8307 11940 8311 11996
rect 8247 11936 8311 11940
rect 8327 11996 8391 12000
rect 8327 11940 8331 11996
rect 8331 11940 8387 11996
rect 8387 11940 8391 11996
rect 8327 11936 8391 11940
rect 8407 11996 8471 12000
rect 8407 11940 8411 11996
rect 8411 11940 8467 11996
rect 8467 11940 8471 11996
rect 8407 11936 8471 11940
rect 10789 11996 10853 12000
rect 10789 11940 10793 11996
rect 10793 11940 10849 11996
rect 10849 11940 10853 11996
rect 10789 11936 10853 11940
rect 10869 11996 10933 12000
rect 10869 11940 10873 11996
rect 10873 11940 10929 11996
rect 10929 11940 10933 11996
rect 10869 11936 10933 11940
rect 10949 11996 11013 12000
rect 10949 11940 10953 11996
rect 10953 11940 11009 11996
rect 11009 11940 11013 11996
rect 10949 11936 11013 11940
rect 11029 11996 11093 12000
rect 11029 11940 11033 11996
rect 11033 11940 11089 11996
rect 11089 11940 11093 11996
rect 11029 11936 11093 11940
rect 2263 11452 2327 11456
rect 2263 11396 2267 11452
rect 2267 11396 2323 11452
rect 2323 11396 2327 11452
rect 2263 11392 2327 11396
rect 2343 11452 2407 11456
rect 2343 11396 2347 11452
rect 2347 11396 2403 11452
rect 2403 11396 2407 11452
rect 2343 11392 2407 11396
rect 2423 11452 2487 11456
rect 2423 11396 2427 11452
rect 2427 11396 2483 11452
rect 2483 11396 2487 11452
rect 2423 11392 2487 11396
rect 2503 11452 2567 11456
rect 2503 11396 2507 11452
rect 2507 11396 2563 11452
rect 2563 11396 2567 11452
rect 2503 11392 2567 11396
rect 4885 11452 4949 11456
rect 4885 11396 4889 11452
rect 4889 11396 4945 11452
rect 4945 11396 4949 11452
rect 4885 11392 4949 11396
rect 4965 11452 5029 11456
rect 4965 11396 4969 11452
rect 4969 11396 5025 11452
rect 5025 11396 5029 11452
rect 4965 11392 5029 11396
rect 5045 11452 5109 11456
rect 5045 11396 5049 11452
rect 5049 11396 5105 11452
rect 5105 11396 5109 11452
rect 5045 11392 5109 11396
rect 5125 11452 5189 11456
rect 5125 11396 5129 11452
rect 5129 11396 5185 11452
rect 5185 11396 5189 11452
rect 5125 11392 5189 11396
rect 7507 11452 7571 11456
rect 7507 11396 7511 11452
rect 7511 11396 7567 11452
rect 7567 11396 7571 11452
rect 7507 11392 7571 11396
rect 7587 11452 7651 11456
rect 7587 11396 7591 11452
rect 7591 11396 7647 11452
rect 7647 11396 7651 11452
rect 7587 11392 7651 11396
rect 7667 11452 7731 11456
rect 7667 11396 7671 11452
rect 7671 11396 7727 11452
rect 7727 11396 7731 11452
rect 7667 11392 7731 11396
rect 7747 11452 7811 11456
rect 7747 11396 7751 11452
rect 7751 11396 7807 11452
rect 7807 11396 7811 11452
rect 7747 11392 7811 11396
rect 10129 11452 10193 11456
rect 10129 11396 10133 11452
rect 10133 11396 10189 11452
rect 10189 11396 10193 11452
rect 10129 11392 10193 11396
rect 10209 11452 10273 11456
rect 10209 11396 10213 11452
rect 10213 11396 10269 11452
rect 10269 11396 10273 11452
rect 10209 11392 10273 11396
rect 10289 11452 10353 11456
rect 10289 11396 10293 11452
rect 10293 11396 10349 11452
rect 10349 11396 10353 11452
rect 10289 11392 10353 11396
rect 10369 11452 10433 11456
rect 10369 11396 10373 11452
rect 10373 11396 10429 11452
rect 10429 11396 10433 11452
rect 10369 11392 10433 11396
rect 2923 10908 2987 10912
rect 2923 10852 2927 10908
rect 2927 10852 2983 10908
rect 2983 10852 2987 10908
rect 2923 10848 2987 10852
rect 3003 10908 3067 10912
rect 3003 10852 3007 10908
rect 3007 10852 3063 10908
rect 3063 10852 3067 10908
rect 3003 10848 3067 10852
rect 3083 10908 3147 10912
rect 3083 10852 3087 10908
rect 3087 10852 3143 10908
rect 3143 10852 3147 10908
rect 3083 10848 3147 10852
rect 3163 10908 3227 10912
rect 3163 10852 3167 10908
rect 3167 10852 3223 10908
rect 3223 10852 3227 10908
rect 3163 10848 3227 10852
rect 5545 10908 5609 10912
rect 5545 10852 5549 10908
rect 5549 10852 5605 10908
rect 5605 10852 5609 10908
rect 5545 10848 5609 10852
rect 5625 10908 5689 10912
rect 5625 10852 5629 10908
rect 5629 10852 5685 10908
rect 5685 10852 5689 10908
rect 5625 10848 5689 10852
rect 5705 10908 5769 10912
rect 5705 10852 5709 10908
rect 5709 10852 5765 10908
rect 5765 10852 5769 10908
rect 5705 10848 5769 10852
rect 5785 10908 5849 10912
rect 5785 10852 5789 10908
rect 5789 10852 5845 10908
rect 5845 10852 5849 10908
rect 5785 10848 5849 10852
rect 8167 10908 8231 10912
rect 8167 10852 8171 10908
rect 8171 10852 8227 10908
rect 8227 10852 8231 10908
rect 8167 10848 8231 10852
rect 8247 10908 8311 10912
rect 8247 10852 8251 10908
rect 8251 10852 8307 10908
rect 8307 10852 8311 10908
rect 8247 10848 8311 10852
rect 8327 10908 8391 10912
rect 8327 10852 8331 10908
rect 8331 10852 8387 10908
rect 8387 10852 8391 10908
rect 8327 10848 8391 10852
rect 8407 10908 8471 10912
rect 8407 10852 8411 10908
rect 8411 10852 8467 10908
rect 8467 10852 8471 10908
rect 8407 10848 8471 10852
rect 10789 10908 10853 10912
rect 10789 10852 10793 10908
rect 10793 10852 10849 10908
rect 10849 10852 10853 10908
rect 10789 10848 10853 10852
rect 10869 10908 10933 10912
rect 10869 10852 10873 10908
rect 10873 10852 10929 10908
rect 10929 10852 10933 10908
rect 10869 10848 10933 10852
rect 10949 10908 11013 10912
rect 10949 10852 10953 10908
rect 10953 10852 11009 10908
rect 11009 10852 11013 10908
rect 10949 10848 11013 10852
rect 11029 10908 11093 10912
rect 11029 10852 11033 10908
rect 11033 10852 11089 10908
rect 11089 10852 11093 10908
rect 11029 10848 11093 10852
rect 2263 10364 2327 10368
rect 2263 10308 2267 10364
rect 2267 10308 2323 10364
rect 2323 10308 2327 10364
rect 2263 10304 2327 10308
rect 2343 10364 2407 10368
rect 2343 10308 2347 10364
rect 2347 10308 2403 10364
rect 2403 10308 2407 10364
rect 2343 10304 2407 10308
rect 2423 10364 2487 10368
rect 2423 10308 2427 10364
rect 2427 10308 2483 10364
rect 2483 10308 2487 10364
rect 2423 10304 2487 10308
rect 2503 10364 2567 10368
rect 2503 10308 2507 10364
rect 2507 10308 2563 10364
rect 2563 10308 2567 10364
rect 2503 10304 2567 10308
rect 4885 10364 4949 10368
rect 4885 10308 4889 10364
rect 4889 10308 4945 10364
rect 4945 10308 4949 10364
rect 4885 10304 4949 10308
rect 4965 10364 5029 10368
rect 4965 10308 4969 10364
rect 4969 10308 5025 10364
rect 5025 10308 5029 10364
rect 4965 10304 5029 10308
rect 5045 10364 5109 10368
rect 5045 10308 5049 10364
rect 5049 10308 5105 10364
rect 5105 10308 5109 10364
rect 5045 10304 5109 10308
rect 5125 10364 5189 10368
rect 5125 10308 5129 10364
rect 5129 10308 5185 10364
rect 5185 10308 5189 10364
rect 5125 10304 5189 10308
rect 7507 10364 7571 10368
rect 7507 10308 7511 10364
rect 7511 10308 7567 10364
rect 7567 10308 7571 10364
rect 7507 10304 7571 10308
rect 7587 10364 7651 10368
rect 7587 10308 7591 10364
rect 7591 10308 7647 10364
rect 7647 10308 7651 10364
rect 7587 10304 7651 10308
rect 7667 10364 7731 10368
rect 7667 10308 7671 10364
rect 7671 10308 7727 10364
rect 7727 10308 7731 10364
rect 7667 10304 7731 10308
rect 7747 10364 7811 10368
rect 7747 10308 7751 10364
rect 7751 10308 7807 10364
rect 7807 10308 7811 10364
rect 7747 10304 7811 10308
rect 10129 10364 10193 10368
rect 10129 10308 10133 10364
rect 10133 10308 10189 10364
rect 10189 10308 10193 10364
rect 10129 10304 10193 10308
rect 10209 10364 10273 10368
rect 10209 10308 10213 10364
rect 10213 10308 10269 10364
rect 10269 10308 10273 10364
rect 10209 10304 10273 10308
rect 10289 10364 10353 10368
rect 10289 10308 10293 10364
rect 10293 10308 10349 10364
rect 10349 10308 10353 10364
rect 10289 10304 10353 10308
rect 10369 10364 10433 10368
rect 10369 10308 10373 10364
rect 10373 10308 10429 10364
rect 10429 10308 10433 10364
rect 10369 10304 10433 10308
rect 2923 9820 2987 9824
rect 2923 9764 2927 9820
rect 2927 9764 2983 9820
rect 2983 9764 2987 9820
rect 2923 9760 2987 9764
rect 3003 9820 3067 9824
rect 3003 9764 3007 9820
rect 3007 9764 3063 9820
rect 3063 9764 3067 9820
rect 3003 9760 3067 9764
rect 3083 9820 3147 9824
rect 3083 9764 3087 9820
rect 3087 9764 3143 9820
rect 3143 9764 3147 9820
rect 3083 9760 3147 9764
rect 3163 9820 3227 9824
rect 3163 9764 3167 9820
rect 3167 9764 3223 9820
rect 3223 9764 3227 9820
rect 3163 9760 3227 9764
rect 5545 9820 5609 9824
rect 5545 9764 5549 9820
rect 5549 9764 5605 9820
rect 5605 9764 5609 9820
rect 5545 9760 5609 9764
rect 5625 9820 5689 9824
rect 5625 9764 5629 9820
rect 5629 9764 5685 9820
rect 5685 9764 5689 9820
rect 5625 9760 5689 9764
rect 5705 9820 5769 9824
rect 5705 9764 5709 9820
rect 5709 9764 5765 9820
rect 5765 9764 5769 9820
rect 5705 9760 5769 9764
rect 5785 9820 5849 9824
rect 5785 9764 5789 9820
rect 5789 9764 5845 9820
rect 5845 9764 5849 9820
rect 5785 9760 5849 9764
rect 8167 9820 8231 9824
rect 8167 9764 8171 9820
rect 8171 9764 8227 9820
rect 8227 9764 8231 9820
rect 8167 9760 8231 9764
rect 8247 9820 8311 9824
rect 8247 9764 8251 9820
rect 8251 9764 8307 9820
rect 8307 9764 8311 9820
rect 8247 9760 8311 9764
rect 8327 9820 8391 9824
rect 8327 9764 8331 9820
rect 8331 9764 8387 9820
rect 8387 9764 8391 9820
rect 8327 9760 8391 9764
rect 8407 9820 8471 9824
rect 8407 9764 8411 9820
rect 8411 9764 8467 9820
rect 8467 9764 8471 9820
rect 8407 9760 8471 9764
rect 10789 9820 10853 9824
rect 10789 9764 10793 9820
rect 10793 9764 10849 9820
rect 10849 9764 10853 9820
rect 10789 9760 10853 9764
rect 10869 9820 10933 9824
rect 10869 9764 10873 9820
rect 10873 9764 10929 9820
rect 10929 9764 10933 9820
rect 10869 9760 10933 9764
rect 10949 9820 11013 9824
rect 10949 9764 10953 9820
rect 10953 9764 11009 9820
rect 11009 9764 11013 9820
rect 10949 9760 11013 9764
rect 11029 9820 11093 9824
rect 11029 9764 11033 9820
rect 11033 9764 11089 9820
rect 11089 9764 11093 9820
rect 11029 9760 11093 9764
rect 2263 9276 2327 9280
rect 2263 9220 2267 9276
rect 2267 9220 2323 9276
rect 2323 9220 2327 9276
rect 2263 9216 2327 9220
rect 2343 9276 2407 9280
rect 2343 9220 2347 9276
rect 2347 9220 2403 9276
rect 2403 9220 2407 9276
rect 2343 9216 2407 9220
rect 2423 9276 2487 9280
rect 2423 9220 2427 9276
rect 2427 9220 2483 9276
rect 2483 9220 2487 9276
rect 2423 9216 2487 9220
rect 2503 9276 2567 9280
rect 2503 9220 2507 9276
rect 2507 9220 2563 9276
rect 2563 9220 2567 9276
rect 2503 9216 2567 9220
rect 4885 9276 4949 9280
rect 4885 9220 4889 9276
rect 4889 9220 4945 9276
rect 4945 9220 4949 9276
rect 4885 9216 4949 9220
rect 4965 9276 5029 9280
rect 4965 9220 4969 9276
rect 4969 9220 5025 9276
rect 5025 9220 5029 9276
rect 4965 9216 5029 9220
rect 5045 9276 5109 9280
rect 5045 9220 5049 9276
rect 5049 9220 5105 9276
rect 5105 9220 5109 9276
rect 5045 9216 5109 9220
rect 5125 9276 5189 9280
rect 5125 9220 5129 9276
rect 5129 9220 5185 9276
rect 5185 9220 5189 9276
rect 5125 9216 5189 9220
rect 7507 9276 7571 9280
rect 7507 9220 7511 9276
rect 7511 9220 7567 9276
rect 7567 9220 7571 9276
rect 7507 9216 7571 9220
rect 7587 9276 7651 9280
rect 7587 9220 7591 9276
rect 7591 9220 7647 9276
rect 7647 9220 7651 9276
rect 7587 9216 7651 9220
rect 7667 9276 7731 9280
rect 7667 9220 7671 9276
rect 7671 9220 7727 9276
rect 7727 9220 7731 9276
rect 7667 9216 7731 9220
rect 7747 9276 7811 9280
rect 7747 9220 7751 9276
rect 7751 9220 7807 9276
rect 7807 9220 7811 9276
rect 7747 9216 7811 9220
rect 10129 9276 10193 9280
rect 10129 9220 10133 9276
rect 10133 9220 10189 9276
rect 10189 9220 10193 9276
rect 10129 9216 10193 9220
rect 10209 9276 10273 9280
rect 10209 9220 10213 9276
rect 10213 9220 10269 9276
rect 10269 9220 10273 9276
rect 10209 9216 10273 9220
rect 10289 9276 10353 9280
rect 10289 9220 10293 9276
rect 10293 9220 10349 9276
rect 10349 9220 10353 9276
rect 10289 9216 10353 9220
rect 10369 9276 10433 9280
rect 10369 9220 10373 9276
rect 10373 9220 10429 9276
rect 10429 9220 10433 9276
rect 10369 9216 10433 9220
rect 2923 8732 2987 8736
rect 2923 8676 2927 8732
rect 2927 8676 2983 8732
rect 2983 8676 2987 8732
rect 2923 8672 2987 8676
rect 3003 8732 3067 8736
rect 3003 8676 3007 8732
rect 3007 8676 3063 8732
rect 3063 8676 3067 8732
rect 3003 8672 3067 8676
rect 3083 8732 3147 8736
rect 3083 8676 3087 8732
rect 3087 8676 3143 8732
rect 3143 8676 3147 8732
rect 3083 8672 3147 8676
rect 3163 8732 3227 8736
rect 3163 8676 3167 8732
rect 3167 8676 3223 8732
rect 3223 8676 3227 8732
rect 3163 8672 3227 8676
rect 5545 8732 5609 8736
rect 5545 8676 5549 8732
rect 5549 8676 5605 8732
rect 5605 8676 5609 8732
rect 5545 8672 5609 8676
rect 5625 8732 5689 8736
rect 5625 8676 5629 8732
rect 5629 8676 5685 8732
rect 5685 8676 5689 8732
rect 5625 8672 5689 8676
rect 5705 8732 5769 8736
rect 5705 8676 5709 8732
rect 5709 8676 5765 8732
rect 5765 8676 5769 8732
rect 5705 8672 5769 8676
rect 5785 8732 5849 8736
rect 5785 8676 5789 8732
rect 5789 8676 5845 8732
rect 5845 8676 5849 8732
rect 5785 8672 5849 8676
rect 8167 8732 8231 8736
rect 8167 8676 8171 8732
rect 8171 8676 8227 8732
rect 8227 8676 8231 8732
rect 8167 8672 8231 8676
rect 8247 8732 8311 8736
rect 8247 8676 8251 8732
rect 8251 8676 8307 8732
rect 8307 8676 8311 8732
rect 8247 8672 8311 8676
rect 8327 8732 8391 8736
rect 8327 8676 8331 8732
rect 8331 8676 8387 8732
rect 8387 8676 8391 8732
rect 8327 8672 8391 8676
rect 8407 8732 8471 8736
rect 8407 8676 8411 8732
rect 8411 8676 8467 8732
rect 8467 8676 8471 8732
rect 8407 8672 8471 8676
rect 10789 8732 10853 8736
rect 10789 8676 10793 8732
rect 10793 8676 10849 8732
rect 10849 8676 10853 8732
rect 10789 8672 10853 8676
rect 10869 8732 10933 8736
rect 10869 8676 10873 8732
rect 10873 8676 10929 8732
rect 10929 8676 10933 8732
rect 10869 8672 10933 8676
rect 10949 8732 11013 8736
rect 10949 8676 10953 8732
rect 10953 8676 11009 8732
rect 11009 8676 11013 8732
rect 10949 8672 11013 8676
rect 11029 8732 11093 8736
rect 11029 8676 11033 8732
rect 11033 8676 11089 8732
rect 11089 8676 11093 8732
rect 11029 8672 11093 8676
rect 2263 8188 2327 8192
rect 2263 8132 2267 8188
rect 2267 8132 2323 8188
rect 2323 8132 2327 8188
rect 2263 8128 2327 8132
rect 2343 8188 2407 8192
rect 2343 8132 2347 8188
rect 2347 8132 2403 8188
rect 2403 8132 2407 8188
rect 2343 8128 2407 8132
rect 2423 8188 2487 8192
rect 2423 8132 2427 8188
rect 2427 8132 2483 8188
rect 2483 8132 2487 8188
rect 2423 8128 2487 8132
rect 2503 8188 2567 8192
rect 2503 8132 2507 8188
rect 2507 8132 2563 8188
rect 2563 8132 2567 8188
rect 2503 8128 2567 8132
rect 4885 8188 4949 8192
rect 4885 8132 4889 8188
rect 4889 8132 4945 8188
rect 4945 8132 4949 8188
rect 4885 8128 4949 8132
rect 4965 8188 5029 8192
rect 4965 8132 4969 8188
rect 4969 8132 5025 8188
rect 5025 8132 5029 8188
rect 4965 8128 5029 8132
rect 5045 8188 5109 8192
rect 5045 8132 5049 8188
rect 5049 8132 5105 8188
rect 5105 8132 5109 8188
rect 5045 8128 5109 8132
rect 5125 8188 5189 8192
rect 5125 8132 5129 8188
rect 5129 8132 5185 8188
rect 5185 8132 5189 8188
rect 5125 8128 5189 8132
rect 7507 8188 7571 8192
rect 7507 8132 7511 8188
rect 7511 8132 7567 8188
rect 7567 8132 7571 8188
rect 7507 8128 7571 8132
rect 7587 8188 7651 8192
rect 7587 8132 7591 8188
rect 7591 8132 7647 8188
rect 7647 8132 7651 8188
rect 7587 8128 7651 8132
rect 7667 8188 7731 8192
rect 7667 8132 7671 8188
rect 7671 8132 7727 8188
rect 7727 8132 7731 8188
rect 7667 8128 7731 8132
rect 7747 8188 7811 8192
rect 7747 8132 7751 8188
rect 7751 8132 7807 8188
rect 7807 8132 7811 8188
rect 7747 8128 7811 8132
rect 10129 8188 10193 8192
rect 10129 8132 10133 8188
rect 10133 8132 10189 8188
rect 10189 8132 10193 8188
rect 10129 8128 10193 8132
rect 10209 8188 10273 8192
rect 10209 8132 10213 8188
rect 10213 8132 10269 8188
rect 10269 8132 10273 8188
rect 10209 8128 10273 8132
rect 10289 8188 10353 8192
rect 10289 8132 10293 8188
rect 10293 8132 10349 8188
rect 10349 8132 10353 8188
rect 10289 8128 10353 8132
rect 10369 8188 10433 8192
rect 10369 8132 10373 8188
rect 10373 8132 10429 8188
rect 10429 8132 10433 8188
rect 10369 8128 10433 8132
rect 2923 7644 2987 7648
rect 2923 7588 2927 7644
rect 2927 7588 2983 7644
rect 2983 7588 2987 7644
rect 2923 7584 2987 7588
rect 3003 7644 3067 7648
rect 3003 7588 3007 7644
rect 3007 7588 3063 7644
rect 3063 7588 3067 7644
rect 3003 7584 3067 7588
rect 3083 7644 3147 7648
rect 3083 7588 3087 7644
rect 3087 7588 3143 7644
rect 3143 7588 3147 7644
rect 3083 7584 3147 7588
rect 3163 7644 3227 7648
rect 3163 7588 3167 7644
rect 3167 7588 3223 7644
rect 3223 7588 3227 7644
rect 3163 7584 3227 7588
rect 5545 7644 5609 7648
rect 5545 7588 5549 7644
rect 5549 7588 5605 7644
rect 5605 7588 5609 7644
rect 5545 7584 5609 7588
rect 5625 7644 5689 7648
rect 5625 7588 5629 7644
rect 5629 7588 5685 7644
rect 5685 7588 5689 7644
rect 5625 7584 5689 7588
rect 5705 7644 5769 7648
rect 5705 7588 5709 7644
rect 5709 7588 5765 7644
rect 5765 7588 5769 7644
rect 5705 7584 5769 7588
rect 5785 7644 5849 7648
rect 5785 7588 5789 7644
rect 5789 7588 5845 7644
rect 5845 7588 5849 7644
rect 5785 7584 5849 7588
rect 8167 7644 8231 7648
rect 8167 7588 8171 7644
rect 8171 7588 8227 7644
rect 8227 7588 8231 7644
rect 8167 7584 8231 7588
rect 8247 7644 8311 7648
rect 8247 7588 8251 7644
rect 8251 7588 8307 7644
rect 8307 7588 8311 7644
rect 8247 7584 8311 7588
rect 8327 7644 8391 7648
rect 8327 7588 8331 7644
rect 8331 7588 8387 7644
rect 8387 7588 8391 7644
rect 8327 7584 8391 7588
rect 8407 7644 8471 7648
rect 8407 7588 8411 7644
rect 8411 7588 8467 7644
rect 8467 7588 8471 7644
rect 8407 7584 8471 7588
rect 10789 7644 10853 7648
rect 10789 7588 10793 7644
rect 10793 7588 10849 7644
rect 10849 7588 10853 7644
rect 10789 7584 10853 7588
rect 10869 7644 10933 7648
rect 10869 7588 10873 7644
rect 10873 7588 10929 7644
rect 10929 7588 10933 7644
rect 10869 7584 10933 7588
rect 10949 7644 11013 7648
rect 10949 7588 10953 7644
rect 10953 7588 11009 7644
rect 11009 7588 11013 7644
rect 10949 7584 11013 7588
rect 11029 7644 11093 7648
rect 11029 7588 11033 7644
rect 11033 7588 11089 7644
rect 11089 7588 11093 7644
rect 11029 7584 11093 7588
rect 2263 7100 2327 7104
rect 2263 7044 2267 7100
rect 2267 7044 2323 7100
rect 2323 7044 2327 7100
rect 2263 7040 2327 7044
rect 2343 7100 2407 7104
rect 2343 7044 2347 7100
rect 2347 7044 2403 7100
rect 2403 7044 2407 7100
rect 2343 7040 2407 7044
rect 2423 7100 2487 7104
rect 2423 7044 2427 7100
rect 2427 7044 2483 7100
rect 2483 7044 2487 7100
rect 2423 7040 2487 7044
rect 2503 7100 2567 7104
rect 2503 7044 2507 7100
rect 2507 7044 2563 7100
rect 2563 7044 2567 7100
rect 2503 7040 2567 7044
rect 4885 7100 4949 7104
rect 4885 7044 4889 7100
rect 4889 7044 4945 7100
rect 4945 7044 4949 7100
rect 4885 7040 4949 7044
rect 4965 7100 5029 7104
rect 4965 7044 4969 7100
rect 4969 7044 5025 7100
rect 5025 7044 5029 7100
rect 4965 7040 5029 7044
rect 5045 7100 5109 7104
rect 5045 7044 5049 7100
rect 5049 7044 5105 7100
rect 5105 7044 5109 7100
rect 5045 7040 5109 7044
rect 5125 7100 5189 7104
rect 5125 7044 5129 7100
rect 5129 7044 5185 7100
rect 5185 7044 5189 7100
rect 5125 7040 5189 7044
rect 7507 7100 7571 7104
rect 7507 7044 7511 7100
rect 7511 7044 7567 7100
rect 7567 7044 7571 7100
rect 7507 7040 7571 7044
rect 7587 7100 7651 7104
rect 7587 7044 7591 7100
rect 7591 7044 7647 7100
rect 7647 7044 7651 7100
rect 7587 7040 7651 7044
rect 7667 7100 7731 7104
rect 7667 7044 7671 7100
rect 7671 7044 7727 7100
rect 7727 7044 7731 7100
rect 7667 7040 7731 7044
rect 7747 7100 7811 7104
rect 7747 7044 7751 7100
rect 7751 7044 7807 7100
rect 7807 7044 7811 7100
rect 7747 7040 7811 7044
rect 10129 7100 10193 7104
rect 10129 7044 10133 7100
rect 10133 7044 10189 7100
rect 10189 7044 10193 7100
rect 10129 7040 10193 7044
rect 10209 7100 10273 7104
rect 10209 7044 10213 7100
rect 10213 7044 10269 7100
rect 10269 7044 10273 7100
rect 10209 7040 10273 7044
rect 10289 7100 10353 7104
rect 10289 7044 10293 7100
rect 10293 7044 10349 7100
rect 10349 7044 10353 7100
rect 10289 7040 10353 7044
rect 10369 7100 10433 7104
rect 10369 7044 10373 7100
rect 10373 7044 10429 7100
rect 10429 7044 10433 7100
rect 10369 7040 10433 7044
rect 2923 6556 2987 6560
rect 2923 6500 2927 6556
rect 2927 6500 2983 6556
rect 2983 6500 2987 6556
rect 2923 6496 2987 6500
rect 3003 6556 3067 6560
rect 3003 6500 3007 6556
rect 3007 6500 3063 6556
rect 3063 6500 3067 6556
rect 3003 6496 3067 6500
rect 3083 6556 3147 6560
rect 3083 6500 3087 6556
rect 3087 6500 3143 6556
rect 3143 6500 3147 6556
rect 3083 6496 3147 6500
rect 3163 6556 3227 6560
rect 3163 6500 3167 6556
rect 3167 6500 3223 6556
rect 3223 6500 3227 6556
rect 3163 6496 3227 6500
rect 5545 6556 5609 6560
rect 5545 6500 5549 6556
rect 5549 6500 5605 6556
rect 5605 6500 5609 6556
rect 5545 6496 5609 6500
rect 5625 6556 5689 6560
rect 5625 6500 5629 6556
rect 5629 6500 5685 6556
rect 5685 6500 5689 6556
rect 5625 6496 5689 6500
rect 5705 6556 5769 6560
rect 5705 6500 5709 6556
rect 5709 6500 5765 6556
rect 5765 6500 5769 6556
rect 5705 6496 5769 6500
rect 5785 6556 5849 6560
rect 5785 6500 5789 6556
rect 5789 6500 5845 6556
rect 5845 6500 5849 6556
rect 5785 6496 5849 6500
rect 8167 6556 8231 6560
rect 8167 6500 8171 6556
rect 8171 6500 8227 6556
rect 8227 6500 8231 6556
rect 8167 6496 8231 6500
rect 8247 6556 8311 6560
rect 8247 6500 8251 6556
rect 8251 6500 8307 6556
rect 8307 6500 8311 6556
rect 8247 6496 8311 6500
rect 8327 6556 8391 6560
rect 8327 6500 8331 6556
rect 8331 6500 8387 6556
rect 8387 6500 8391 6556
rect 8327 6496 8391 6500
rect 8407 6556 8471 6560
rect 8407 6500 8411 6556
rect 8411 6500 8467 6556
rect 8467 6500 8471 6556
rect 8407 6496 8471 6500
rect 10789 6556 10853 6560
rect 10789 6500 10793 6556
rect 10793 6500 10849 6556
rect 10849 6500 10853 6556
rect 10789 6496 10853 6500
rect 10869 6556 10933 6560
rect 10869 6500 10873 6556
rect 10873 6500 10929 6556
rect 10929 6500 10933 6556
rect 10869 6496 10933 6500
rect 10949 6556 11013 6560
rect 10949 6500 10953 6556
rect 10953 6500 11009 6556
rect 11009 6500 11013 6556
rect 10949 6496 11013 6500
rect 11029 6556 11093 6560
rect 11029 6500 11033 6556
rect 11033 6500 11089 6556
rect 11089 6500 11093 6556
rect 11029 6496 11093 6500
rect 2263 6012 2327 6016
rect 2263 5956 2267 6012
rect 2267 5956 2323 6012
rect 2323 5956 2327 6012
rect 2263 5952 2327 5956
rect 2343 6012 2407 6016
rect 2343 5956 2347 6012
rect 2347 5956 2403 6012
rect 2403 5956 2407 6012
rect 2343 5952 2407 5956
rect 2423 6012 2487 6016
rect 2423 5956 2427 6012
rect 2427 5956 2483 6012
rect 2483 5956 2487 6012
rect 2423 5952 2487 5956
rect 2503 6012 2567 6016
rect 2503 5956 2507 6012
rect 2507 5956 2563 6012
rect 2563 5956 2567 6012
rect 2503 5952 2567 5956
rect 4885 6012 4949 6016
rect 4885 5956 4889 6012
rect 4889 5956 4945 6012
rect 4945 5956 4949 6012
rect 4885 5952 4949 5956
rect 4965 6012 5029 6016
rect 4965 5956 4969 6012
rect 4969 5956 5025 6012
rect 5025 5956 5029 6012
rect 4965 5952 5029 5956
rect 5045 6012 5109 6016
rect 5045 5956 5049 6012
rect 5049 5956 5105 6012
rect 5105 5956 5109 6012
rect 5045 5952 5109 5956
rect 5125 6012 5189 6016
rect 5125 5956 5129 6012
rect 5129 5956 5185 6012
rect 5185 5956 5189 6012
rect 5125 5952 5189 5956
rect 7507 6012 7571 6016
rect 7507 5956 7511 6012
rect 7511 5956 7567 6012
rect 7567 5956 7571 6012
rect 7507 5952 7571 5956
rect 7587 6012 7651 6016
rect 7587 5956 7591 6012
rect 7591 5956 7647 6012
rect 7647 5956 7651 6012
rect 7587 5952 7651 5956
rect 7667 6012 7731 6016
rect 7667 5956 7671 6012
rect 7671 5956 7727 6012
rect 7727 5956 7731 6012
rect 7667 5952 7731 5956
rect 7747 6012 7811 6016
rect 7747 5956 7751 6012
rect 7751 5956 7807 6012
rect 7807 5956 7811 6012
rect 7747 5952 7811 5956
rect 10129 6012 10193 6016
rect 10129 5956 10133 6012
rect 10133 5956 10189 6012
rect 10189 5956 10193 6012
rect 10129 5952 10193 5956
rect 10209 6012 10273 6016
rect 10209 5956 10213 6012
rect 10213 5956 10269 6012
rect 10269 5956 10273 6012
rect 10209 5952 10273 5956
rect 10289 6012 10353 6016
rect 10289 5956 10293 6012
rect 10293 5956 10349 6012
rect 10349 5956 10353 6012
rect 10289 5952 10353 5956
rect 10369 6012 10433 6016
rect 10369 5956 10373 6012
rect 10373 5956 10429 6012
rect 10429 5956 10433 6012
rect 10369 5952 10433 5956
rect 2923 5468 2987 5472
rect 2923 5412 2927 5468
rect 2927 5412 2983 5468
rect 2983 5412 2987 5468
rect 2923 5408 2987 5412
rect 3003 5468 3067 5472
rect 3003 5412 3007 5468
rect 3007 5412 3063 5468
rect 3063 5412 3067 5468
rect 3003 5408 3067 5412
rect 3083 5468 3147 5472
rect 3083 5412 3087 5468
rect 3087 5412 3143 5468
rect 3143 5412 3147 5468
rect 3083 5408 3147 5412
rect 3163 5468 3227 5472
rect 3163 5412 3167 5468
rect 3167 5412 3223 5468
rect 3223 5412 3227 5468
rect 3163 5408 3227 5412
rect 5545 5468 5609 5472
rect 5545 5412 5549 5468
rect 5549 5412 5605 5468
rect 5605 5412 5609 5468
rect 5545 5408 5609 5412
rect 5625 5468 5689 5472
rect 5625 5412 5629 5468
rect 5629 5412 5685 5468
rect 5685 5412 5689 5468
rect 5625 5408 5689 5412
rect 5705 5468 5769 5472
rect 5705 5412 5709 5468
rect 5709 5412 5765 5468
rect 5765 5412 5769 5468
rect 5705 5408 5769 5412
rect 5785 5468 5849 5472
rect 5785 5412 5789 5468
rect 5789 5412 5845 5468
rect 5845 5412 5849 5468
rect 5785 5408 5849 5412
rect 8167 5468 8231 5472
rect 8167 5412 8171 5468
rect 8171 5412 8227 5468
rect 8227 5412 8231 5468
rect 8167 5408 8231 5412
rect 8247 5468 8311 5472
rect 8247 5412 8251 5468
rect 8251 5412 8307 5468
rect 8307 5412 8311 5468
rect 8247 5408 8311 5412
rect 8327 5468 8391 5472
rect 8327 5412 8331 5468
rect 8331 5412 8387 5468
rect 8387 5412 8391 5468
rect 8327 5408 8391 5412
rect 8407 5468 8471 5472
rect 8407 5412 8411 5468
rect 8411 5412 8467 5468
rect 8467 5412 8471 5468
rect 8407 5408 8471 5412
rect 10789 5468 10853 5472
rect 10789 5412 10793 5468
rect 10793 5412 10849 5468
rect 10849 5412 10853 5468
rect 10789 5408 10853 5412
rect 10869 5468 10933 5472
rect 10869 5412 10873 5468
rect 10873 5412 10929 5468
rect 10929 5412 10933 5468
rect 10869 5408 10933 5412
rect 10949 5468 11013 5472
rect 10949 5412 10953 5468
rect 10953 5412 11009 5468
rect 11009 5412 11013 5468
rect 10949 5408 11013 5412
rect 11029 5468 11093 5472
rect 11029 5412 11033 5468
rect 11033 5412 11089 5468
rect 11089 5412 11093 5468
rect 11029 5408 11093 5412
rect 2263 4924 2327 4928
rect 2263 4868 2267 4924
rect 2267 4868 2323 4924
rect 2323 4868 2327 4924
rect 2263 4864 2327 4868
rect 2343 4924 2407 4928
rect 2343 4868 2347 4924
rect 2347 4868 2403 4924
rect 2403 4868 2407 4924
rect 2343 4864 2407 4868
rect 2423 4924 2487 4928
rect 2423 4868 2427 4924
rect 2427 4868 2483 4924
rect 2483 4868 2487 4924
rect 2423 4864 2487 4868
rect 2503 4924 2567 4928
rect 2503 4868 2507 4924
rect 2507 4868 2563 4924
rect 2563 4868 2567 4924
rect 2503 4864 2567 4868
rect 4885 4924 4949 4928
rect 4885 4868 4889 4924
rect 4889 4868 4945 4924
rect 4945 4868 4949 4924
rect 4885 4864 4949 4868
rect 4965 4924 5029 4928
rect 4965 4868 4969 4924
rect 4969 4868 5025 4924
rect 5025 4868 5029 4924
rect 4965 4864 5029 4868
rect 5045 4924 5109 4928
rect 5045 4868 5049 4924
rect 5049 4868 5105 4924
rect 5105 4868 5109 4924
rect 5045 4864 5109 4868
rect 5125 4924 5189 4928
rect 5125 4868 5129 4924
rect 5129 4868 5185 4924
rect 5185 4868 5189 4924
rect 5125 4864 5189 4868
rect 7507 4924 7571 4928
rect 7507 4868 7511 4924
rect 7511 4868 7567 4924
rect 7567 4868 7571 4924
rect 7507 4864 7571 4868
rect 7587 4924 7651 4928
rect 7587 4868 7591 4924
rect 7591 4868 7647 4924
rect 7647 4868 7651 4924
rect 7587 4864 7651 4868
rect 7667 4924 7731 4928
rect 7667 4868 7671 4924
rect 7671 4868 7727 4924
rect 7727 4868 7731 4924
rect 7667 4864 7731 4868
rect 7747 4924 7811 4928
rect 7747 4868 7751 4924
rect 7751 4868 7807 4924
rect 7807 4868 7811 4924
rect 7747 4864 7811 4868
rect 10129 4924 10193 4928
rect 10129 4868 10133 4924
rect 10133 4868 10189 4924
rect 10189 4868 10193 4924
rect 10129 4864 10193 4868
rect 10209 4924 10273 4928
rect 10209 4868 10213 4924
rect 10213 4868 10269 4924
rect 10269 4868 10273 4924
rect 10209 4864 10273 4868
rect 10289 4924 10353 4928
rect 10289 4868 10293 4924
rect 10293 4868 10349 4924
rect 10349 4868 10353 4924
rect 10289 4864 10353 4868
rect 10369 4924 10433 4928
rect 10369 4868 10373 4924
rect 10373 4868 10429 4924
rect 10429 4868 10433 4924
rect 10369 4864 10433 4868
rect 2923 4380 2987 4384
rect 2923 4324 2927 4380
rect 2927 4324 2983 4380
rect 2983 4324 2987 4380
rect 2923 4320 2987 4324
rect 3003 4380 3067 4384
rect 3003 4324 3007 4380
rect 3007 4324 3063 4380
rect 3063 4324 3067 4380
rect 3003 4320 3067 4324
rect 3083 4380 3147 4384
rect 3083 4324 3087 4380
rect 3087 4324 3143 4380
rect 3143 4324 3147 4380
rect 3083 4320 3147 4324
rect 3163 4380 3227 4384
rect 3163 4324 3167 4380
rect 3167 4324 3223 4380
rect 3223 4324 3227 4380
rect 3163 4320 3227 4324
rect 5545 4380 5609 4384
rect 5545 4324 5549 4380
rect 5549 4324 5605 4380
rect 5605 4324 5609 4380
rect 5545 4320 5609 4324
rect 5625 4380 5689 4384
rect 5625 4324 5629 4380
rect 5629 4324 5685 4380
rect 5685 4324 5689 4380
rect 5625 4320 5689 4324
rect 5705 4380 5769 4384
rect 5705 4324 5709 4380
rect 5709 4324 5765 4380
rect 5765 4324 5769 4380
rect 5705 4320 5769 4324
rect 5785 4380 5849 4384
rect 5785 4324 5789 4380
rect 5789 4324 5845 4380
rect 5845 4324 5849 4380
rect 5785 4320 5849 4324
rect 8167 4380 8231 4384
rect 8167 4324 8171 4380
rect 8171 4324 8227 4380
rect 8227 4324 8231 4380
rect 8167 4320 8231 4324
rect 8247 4380 8311 4384
rect 8247 4324 8251 4380
rect 8251 4324 8307 4380
rect 8307 4324 8311 4380
rect 8247 4320 8311 4324
rect 8327 4380 8391 4384
rect 8327 4324 8331 4380
rect 8331 4324 8387 4380
rect 8387 4324 8391 4380
rect 8327 4320 8391 4324
rect 8407 4380 8471 4384
rect 8407 4324 8411 4380
rect 8411 4324 8467 4380
rect 8467 4324 8471 4380
rect 8407 4320 8471 4324
rect 10789 4380 10853 4384
rect 10789 4324 10793 4380
rect 10793 4324 10849 4380
rect 10849 4324 10853 4380
rect 10789 4320 10853 4324
rect 10869 4380 10933 4384
rect 10869 4324 10873 4380
rect 10873 4324 10929 4380
rect 10929 4324 10933 4380
rect 10869 4320 10933 4324
rect 10949 4380 11013 4384
rect 10949 4324 10953 4380
rect 10953 4324 11009 4380
rect 11009 4324 11013 4380
rect 10949 4320 11013 4324
rect 11029 4380 11093 4384
rect 11029 4324 11033 4380
rect 11033 4324 11089 4380
rect 11089 4324 11093 4380
rect 11029 4320 11093 4324
rect 2263 3836 2327 3840
rect 2263 3780 2267 3836
rect 2267 3780 2323 3836
rect 2323 3780 2327 3836
rect 2263 3776 2327 3780
rect 2343 3836 2407 3840
rect 2343 3780 2347 3836
rect 2347 3780 2403 3836
rect 2403 3780 2407 3836
rect 2343 3776 2407 3780
rect 2423 3836 2487 3840
rect 2423 3780 2427 3836
rect 2427 3780 2483 3836
rect 2483 3780 2487 3836
rect 2423 3776 2487 3780
rect 2503 3836 2567 3840
rect 2503 3780 2507 3836
rect 2507 3780 2563 3836
rect 2563 3780 2567 3836
rect 2503 3776 2567 3780
rect 4885 3836 4949 3840
rect 4885 3780 4889 3836
rect 4889 3780 4945 3836
rect 4945 3780 4949 3836
rect 4885 3776 4949 3780
rect 4965 3836 5029 3840
rect 4965 3780 4969 3836
rect 4969 3780 5025 3836
rect 5025 3780 5029 3836
rect 4965 3776 5029 3780
rect 5045 3836 5109 3840
rect 5045 3780 5049 3836
rect 5049 3780 5105 3836
rect 5105 3780 5109 3836
rect 5045 3776 5109 3780
rect 5125 3836 5189 3840
rect 5125 3780 5129 3836
rect 5129 3780 5185 3836
rect 5185 3780 5189 3836
rect 5125 3776 5189 3780
rect 7507 3836 7571 3840
rect 7507 3780 7511 3836
rect 7511 3780 7567 3836
rect 7567 3780 7571 3836
rect 7507 3776 7571 3780
rect 7587 3836 7651 3840
rect 7587 3780 7591 3836
rect 7591 3780 7647 3836
rect 7647 3780 7651 3836
rect 7587 3776 7651 3780
rect 7667 3836 7731 3840
rect 7667 3780 7671 3836
rect 7671 3780 7727 3836
rect 7727 3780 7731 3836
rect 7667 3776 7731 3780
rect 7747 3836 7811 3840
rect 7747 3780 7751 3836
rect 7751 3780 7807 3836
rect 7807 3780 7811 3836
rect 7747 3776 7811 3780
rect 10129 3836 10193 3840
rect 10129 3780 10133 3836
rect 10133 3780 10189 3836
rect 10189 3780 10193 3836
rect 10129 3776 10193 3780
rect 10209 3836 10273 3840
rect 10209 3780 10213 3836
rect 10213 3780 10269 3836
rect 10269 3780 10273 3836
rect 10209 3776 10273 3780
rect 10289 3836 10353 3840
rect 10289 3780 10293 3836
rect 10293 3780 10349 3836
rect 10349 3780 10353 3836
rect 10289 3776 10353 3780
rect 10369 3836 10433 3840
rect 10369 3780 10373 3836
rect 10373 3780 10429 3836
rect 10429 3780 10433 3836
rect 10369 3776 10433 3780
rect 2923 3292 2987 3296
rect 2923 3236 2927 3292
rect 2927 3236 2983 3292
rect 2983 3236 2987 3292
rect 2923 3232 2987 3236
rect 3003 3292 3067 3296
rect 3003 3236 3007 3292
rect 3007 3236 3063 3292
rect 3063 3236 3067 3292
rect 3003 3232 3067 3236
rect 3083 3292 3147 3296
rect 3083 3236 3087 3292
rect 3087 3236 3143 3292
rect 3143 3236 3147 3292
rect 3083 3232 3147 3236
rect 3163 3292 3227 3296
rect 3163 3236 3167 3292
rect 3167 3236 3223 3292
rect 3223 3236 3227 3292
rect 3163 3232 3227 3236
rect 5545 3292 5609 3296
rect 5545 3236 5549 3292
rect 5549 3236 5605 3292
rect 5605 3236 5609 3292
rect 5545 3232 5609 3236
rect 5625 3292 5689 3296
rect 5625 3236 5629 3292
rect 5629 3236 5685 3292
rect 5685 3236 5689 3292
rect 5625 3232 5689 3236
rect 5705 3292 5769 3296
rect 5705 3236 5709 3292
rect 5709 3236 5765 3292
rect 5765 3236 5769 3292
rect 5705 3232 5769 3236
rect 5785 3292 5849 3296
rect 5785 3236 5789 3292
rect 5789 3236 5845 3292
rect 5845 3236 5849 3292
rect 5785 3232 5849 3236
rect 8167 3292 8231 3296
rect 8167 3236 8171 3292
rect 8171 3236 8227 3292
rect 8227 3236 8231 3292
rect 8167 3232 8231 3236
rect 8247 3292 8311 3296
rect 8247 3236 8251 3292
rect 8251 3236 8307 3292
rect 8307 3236 8311 3292
rect 8247 3232 8311 3236
rect 8327 3292 8391 3296
rect 8327 3236 8331 3292
rect 8331 3236 8387 3292
rect 8387 3236 8391 3292
rect 8327 3232 8391 3236
rect 8407 3292 8471 3296
rect 8407 3236 8411 3292
rect 8411 3236 8467 3292
rect 8467 3236 8471 3292
rect 8407 3232 8471 3236
rect 10789 3292 10853 3296
rect 10789 3236 10793 3292
rect 10793 3236 10849 3292
rect 10849 3236 10853 3292
rect 10789 3232 10853 3236
rect 10869 3292 10933 3296
rect 10869 3236 10873 3292
rect 10873 3236 10929 3292
rect 10929 3236 10933 3292
rect 10869 3232 10933 3236
rect 10949 3292 11013 3296
rect 10949 3236 10953 3292
rect 10953 3236 11009 3292
rect 11009 3236 11013 3292
rect 10949 3232 11013 3236
rect 11029 3292 11093 3296
rect 11029 3236 11033 3292
rect 11033 3236 11089 3292
rect 11089 3236 11093 3292
rect 11029 3232 11093 3236
rect 2263 2748 2327 2752
rect 2263 2692 2267 2748
rect 2267 2692 2323 2748
rect 2323 2692 2327 2748
rect 2263 2688 2327 2692
rect 2343 2748 2407 2752
rect 2343 2692 2347 2748
rect 2347 2692 2403 2748
rect 2403 2692 2407 2748
rect 2343 2688 2407 2692
rect 2423 2748 2487 2752
rect 2423 2692 2427 2748
rect 2427 2692 2483 2748
rect 2483 2692 2487 2748
rect 2423 2688 2487 2692
rect 2503 2748 2567 2752
rect 2503 2692 2507 2748
rect 2507 2692 2563 2748
rect 2563 2692 2567 2748
rect 2503 2688 2567 2692
rect 4885 2748 4949 2752
rect 4885 2692 4889 2748
rect 4889 2692 4945 2748
rect 4945 2692 4949 2748
rect 4885 2688 4949 2692
rect 4965 2748 5029 2752
rect 4965 2692 4969 2748
rect 4969 2692 5025 2748
rect 5025 2692 5029 2748
rect 4965 2688 5029 2692
rect 5045 2748 5109 2752
rect 5045 2692 5049 2748
rect 5049 2692 5105 2748
rect 5105 2692 5109 2748
rect 5045 2688 5109 2692
rect 5125 2748 5189 2752
rect 5125 2692 5129 2748
rect 5129 2692 5185 2748
rect 5185 2692 5189 2748
rect 5125 2688 5189 2692
rect 7507 2748 7571 2752
rect 7507 2692 7511 2748
rect 7511 2692 7567 2748
rect 7567 2692 7571 2748
rect 7507 2688 7571 2692
rect 7587 2748 7651 2752
rect 7587 2692 7591 2748
rect 7591 2692 7647 2748
rect 7647 2692 7651 2748
rect 7587 2688 7651 2692
rect 7667 2748 7731 2752
rect 7667 2692 7671 2748
rect 7671 2692 7727 2748
rect 7727 2692 7731 2748
rect 7667 2688 7731 2692
rect 7747 2748 7811 2752
rect 7747 2692 7751 2748
rect 7751 2692 7807 2748
rect 7807 2692 7811 2748
rect 7747 2688 7811 2692
rect 10129 2748 10193 2752
rect 10129 2692 10133 2748
rect 10133 2692 10189 2748
rect 10189 2692 10193 2748
rect 10129 2688 10193 2692
rect 10209 2748 10273 2752
rect 10209 2692 10213 2748
rect 10213 2692 10269 2748
rect 10269 2692 10273 2748
rect 10209 2688 10273 2692
rect 10289 2748 10353 2752
rect 10289 2692 10293 2748
rect 10293 2692 10349 2748
rect 10349 2692 10353 2748
rect 10289 2688 10353 2692
rect 10369 2748 10433 2752
rect 10369 2692 10373 2748
rect 10373 2692 10429 2748
rect 10429 2692 10433 2748
rect 10369 2688 10433 2692
rect 2923 2204 2987 2208
rect 2923 2148 2927 2204
rect 2927 2148 2983 2204
rect 2983 2148 2987 2204
rect 2923 2144 2987 2148
rect 3003 2204 3067 2208
rect 3003 2148 3007 2204
rect 3007 2148 3063 2204
rect 3063 2148 3067 2204
rect 3003 2144 3067 2148
rect 3083 2204 3147 2208
rect 3083 2148 3087 2204
rect 3087 2148 3143 2204
rect 3143 2148 3147 2204
rect 3083 2144 3147 2148
rect 3163 2204 3227 2208
rect 3163 2148 3167 2204
rect 3167 2148 3223 2204
rect 3223 2148 3227 2204
rect 3163 2144 3227 2148
rect 5545 2204 5609 2208
rect 5545 2148 5549 2204
rect 5549 2148 5605 2204
rect 5605 2148 5609 2204
rect 5545 2144 5609 2148
rect 5625 2204 5689 2208
rect 5625 2148 5629 2204
rect 5629 2148 5685 2204
rect 5685 2148 5689 2204
rect 5625 2144 5689 2148
rect 5705 2204 5769 2208
rect 5705 2148 5709 2204
rect 5709 2148 5765 2204
rect 5765 2148 5769 2204
rect 5705 2144 5769 2148
rect 5785 2204 5849 2208
rect 5785 2148 5789 2204
rect 5789 2148 5845 2204
rect 5845 2148 5849 2204
rect 5785 2144 5849 2148
rect 8167 2204 8231 2208
rect 8167 2148 8171 2204
rect 8171 2148 8227 2204
rect 8227 2148 8231 2204
rect 8167 2144 8231 2148
rect 8247 2204 8311 2208
rect 8247 2148 8251 2204
rect 8251 2148 8307 2204
rect 8307 2148 8311 2204
rect 8247 2144 8311 2148
rect 8327 2204 8391 2208
rect 8327 2148 8331 2204
rect 8331 2148 8387 2204
rect 8387 2148 8391 2204
rect 8327 2144 8391 2148
rect 8407 2204 8471 2208
rect 8407 2148 8411 2204
rect 8411 2148 8467 2204
rect 8467 2148 8471 2204
rect 8407 2144 8471 2148
rect 10789 2204 10853 2208
rect 10789 2148 10793 2204
rect 10793 2148 10849 2204
rect 10849 2148 10853 2204
rect 10789 2144 10853 2148
rect 10869 2204 10933 2208
rect 10869 2148 10873 2204
rect 10873 2148 10929 2204
rect 10929 2148 10933 2204
rect 10869 2144 10933 2148
rect 10949 2204 11013 2208
rect 10949 2148 10953 2204
rect 10953 2148 11009 2204
rect 11009 2148 11013 2204
rect 10949 2144 11013 2148
rect 11029 2204 11093 2208
rect 11029 2148 11033 2204
rect 11033 2148 11089 2204
rect 11089 2148 11093 2204
rect 11029 2144 11093 2148
<< metal4 >>
rect 2255 12544 2575 12560
rect 2255 12480 2263 12544
rect 2327 12480 2343 12544
rect 2407 12480 2423 12544
rect 2487 12480 2503 12544
rect 2567 12480 2575 12544
rect 2255 11456 2575 12480
rect 2255 11392 2263 11456
rect 2327 11392 2343 11456
rect 2407 11392 2423 11456
rect 2487 11392 2503 11456
rect 2567 11392 2575 11456
rect 2255 11338 2575 11392
rect 2255 11102 2297 11338
rect 2533 11102 2575 11338
rect 2255 10368 2575 11102
rect 2255 10304 2263 10368
rect 2327 10304 2343 10368
rect 2407 10304 2423 10368
rect 2487 10304 2503 10368
rect 2567 10304 2575 10368
rect 2255 9280 2575 10304
rect 2255 9216 2263 9280
rect 2327 9216 2343 9280
rect 2407 9216 2423 9280
rect 2487 9216 2503 9280
rect 2567 9216 2575 9280
rect 2255 8754 2575 9216
rect 2255 8518 2297 8754
rect 2533 8518 2575 8754
rect 2255 8192 2575 8518
rect 2255 8128 2263 8192
rect 2327 8128 2343 8192
rect 2407 8128 2423 8192
rect 2487 8128 2503 8192
rect 2567 8128 2575 8192
rect 2255 7104 2575 8128
rect 2255 7040 2263 7104
rect 2327 7040 2343 7104
rect 2407 7040 2423 7104
rect 2487 7040 2503 7104
rect 2567 7040 2575 7104
rect 2255 6170 2575 7040
rect 2255 6016 2297 6170
rect 2533 6016 2575 6170
rect 2255 5952 2263 6016
rect 2567 5952 2575 6016
rect 2255 5934 2297 5952
rect 2533 5934 2575 5952
rect 2255 4928 2575 5934
rect 2255 4864 2263 4928
rect 2327 4864 2343 4928
rect 2407 4864 2423 4928
rect 2487 4864 2503 4928
rect 2567 4864 2575 4928
rect 2255 3840 2575 4864
rect 2255 3776 2263 3840
rect 2327 3776 2343 3840
rect 2407 3776 2423 3840
rect 2487 3776 2503 3840
rect 2567 3776 2575 3840
rect 2255 3586 2575 3776
rect 2255 3350 2297 3586
rect 2533 3350 2575 3586
rect 2255 2752 2575 3350
rect 2255 2688 2263 2752
rect 2327 2688 2343 2752
rect 2407 2688 2423 2752
rect 2487 2688 2503 2752
rect 2567 2688 2575 2752
rect 2255 2128 2575 2688
rect 2915 12000 3235 12560
rect 2915 11936 2923 12000
rect 2987 11998 3003 12000
rect 3067 11998 3083 12000
rect 3147 11998 3163 12000
rect 3227 11936 3235 12000
rect 2915 11762 2957 11936
rect 3193 11762 3235 11936
rect 2915 10912 3235 11762
rect 2915 10848 2923 10912
rect 2987 10848 3003 10912
rect 3067 10848 3083 10912
rect 3147 10848 3163 10912
rect 3227 10848 3235 10912
rect 2915 9824 3235 10848
rect 2915 9760 2923 9824
rect 2987 9760 3003 9824
rect 3067 9760 3083 9824
rect 3147 9760 3163 9824
rect 3227 9760 3235 9824
rect 2915 9414 3235 9760
rect 2915 9178 2957 9414
rect 3193 9178 3235 9414
rect 2915 8736 3235 9178
rect 2915 8672 2923 8736
rect 2987 8672 3003 8736
rect 3067 8672 3083 8736
rect 3147 8672 3163 8736
rect 3227 8672 3235 8736
rect 2915 7648 3235 8672
rect 2915 7584 2923 7648
rect 2987 7584 3003 7648
rect 3067 7584 3083 7648
rect 3147 7584 3163 7648
rect 3227 7584 3235 7648
rect 2915 6830 3235 7584
rect 2915 6594 2957 6830
rect 3193 6594 3235 6830
rect 2915 6560 3235 6594
rect 2915 6496 2923 6560
rect 2987 6496 3003 6560
rect 3067 6496 3083 6560
rect 3147 6496 3163 6560
rect 3227 6496 3235 6560
rect 2915 5472 3235 6496
rect 2915 5408 2923 5472
rect 2987 5408 3003 5472
rect 3067 5408 3083 5472
rect 3147 5408 3163 5472
rect 3227 5408 3235 5472
rect 2915 4384 3235 5408
rect 2915 4320 2923 4384
rect 2987 4320 3003 4384
rect 3067 4320 3083 4384
rect 3147 4320 3163 4384
rect 3227 4320 3235 4384
rect 2915 4246 3235 4320
rect 2915 4010 2957 4246
rect 3193 4010 3235 4246
rect 2915 3296 3235 4010
rect 2915 3232 2923 3296
rect 2987 3232 3003 3296
rect 3067 3232 3083 3296
rect 3147 3232 3163 3296
rect 3227 3232 3235 3296
rect 2915 2208 3235 3232
rect 2915 2144 2923 2208
rect 2987 2144 3003 2208
rect 3067 2144 3083 2208
rect 3147 2144 3163 2208
rect 3227 2144 3235 2208
rect 2915 2128 3235 2144
rect 4877 12544 5197 12560
rect 4877 12480 4885 12544
rect 4949 12480 4965 12544
rect 5029 12480 5045 12544
rect 5109 12480 5125 12544
rect 5189 12480 5197 12544
rect 4877 11456 5197 12480
rect 4877 11392 4885 11456
rect 4949 11392 4965 11456
rect 5029 11392 5045 11456
rect 5109 11392 5125 11456
rect 5189 11392 5197 11456
rect 4877 11338 5197 11392
rect 4877 11102 4919 11338
rect 5155 11102 5197 11338
rect 4877 10368 5197 11102
rect 4877 10304 4885 10368
rect 4949 10304 4965 10368
rect 5029 10304 5045 10368
rect 5109 10304 5125 10368
rect 5189 10304 5197 10368
rect 4877 9280 5197 10304
rect 4877 9216 4885 9280
rect 4949 9216 4965 9280
rect 5029 9216 5045 9280
rect 5109 9216 5125 9280
rect 5189 9216 5197 9280
rect 4877 8754 5197 9216
rect 4877 8518 4919 8754
rect 5155 8518 5197 8754
rect 4877 8192 5197 8518
rect 4877 8128 4885 8192
rect 4949 8128 4965 8192
rect 5029 8128 5045 8192
rect 5109 8128 5125 8192
rect 5189 8128 5197 8192
rect 4877 7104 5197 8128
rect 4877 7040 4885 7104
rect 4949 7040 4965 7104
rect 5029 7040 5045 7104
rect 5109 7040 5125 7104
rect 5189 7040 5197 7104
rect 4877 6170 5197 7040
rect 4877 6016 4919 6170
rect 5155 6016 5197 6170
rect 4877 5952 4885 6016
rect 5189 5952 5197 6016
rect 4877 5934 4919 5952
rect 5155 5934 5197 5952
rect 4877 4928 5197 5934
rect 4877 4864 4885 4928
rect 4949 4864 4965 4928
rect 5029 4864 5045 4928
rect 5109 4864 5125 4928
rect 5189 4864 5197 4928
rect 4877 3840 5197 4864
rect 4877 3776 4885 3840
rect 4949 3776 4965 3840
rect 5029 3776 5045 3840
rect 5109 3776 5125 3840
rect 5189 3776 5197 3840
rect 4877 3586 5197 3776
rect 4877 3350 4919 3586
rect 5155 3350 5197 3586
rect 4877 2752 5197 3350
rect 4877 2688 4885 2752
rect 4949 2688 4965 2752
rect 5029 2688 5045 2752
rect 5109 2688 5125 2752
rect 5189 2688 5197 2752
rect 4877 2128 5197 2688
rect 5537 12000 5857 12560
rect 5537 11936 5545 12000
rect 5609 11998 5625 12000
rect 5689 11998 5705 12000
rect 5769 11998 5785 12000
rect 5849 11936 5857 12000
rect 5537 11762 5579 11936
rect 5815 11762 5857 11936
rect 5537 10912 5857 11762
rect 5537 10848 5545 10912
rect 5609 10848 5625 10912
rect 5689 10848 5705 10912
rect 5769 10848 5785 10912
rect 5849 10848 5857 10912
rect 5537 9824 5857 10848
rect 5537 9760 5545 9824
rect 5609 9760 5625 9824
rect 5689 9760 5705 9824
rect 5769 9760 5785 9824
rect 5849 9760 5857 9824
rect 5537 9414 5857 9760
rect 5537 9178 5579 9414
rect 5815 9178 5857 9414
rect 5537 8736 5857 9178
rect 5537 8672 5545 8736
rect 5609 8672 5625 8736
rect 5689 8672 5705 8736
rect 5769 8672 5785 8736
rect 5849 8672 5857 8736
rect 5537 7648 5857 8672
rect 5537 7584 5545 7648
rect 5609 7584 5625 7648
rect 5689 7584 5705 7648
rect 5769 7584 5785 7648
rect 5849 7584 5857 7648
rect 5537 6830 5857 7584
rect 5537 6594 5579 6830
rect 5815 6594 5857 6830
rect 5537 6560 5857 6594
rect 5537 6496 5545 6560
rect 5609 6496 5625 6560
rect 5689 6496 5705 6560
rect 5769 6496 5785 6560
rect 5849 6496 5857 6560
rect 5537 5472 5857 6496
rect 5537 5408 5545 5472
rect 5609 5408 5625 5472
rect 5689 5408 5705 5472
rect 5769 5408 5785 5472
rect 5849 5408 5857 5472
rect 5537 4384 5857 5408
rect 5537 4320 5545 4384
rect 5609 4320 5625 4384
rect 5689 4320 5705 4384
rect 5769 4320 5785 4384
rect 5849 4320 5857 4384
rect 5537 4246 5857 4320
rect 5537 4010 5579 4246
rect 5815 4010 5857 4246
rect 5537 3296 5857 4010
rect 5537 3232 5545 3296
rect 5609 3232 5625 3296
rect 5689 3232 5705 3296
rect 5769 3232 5785 3296
rect 5849 3232 5857 3296
rect 5537 2208 5857 3232
rect 5537 2144 5545 2208
rect 5609 2144 5625 2208
rect 5689 2144 5705 2208
rect 5769 2144 5785 2208
rect 5849 2144 5857 2208
rect 5537 2128 5857 2144
rect 7499 12544 7819 12560
rect 7499 12480 7507 12544
rect 7571 12480 7587 12544
rect 7651 12480 7667 12544
rect 7731 12480 7747 12544
rect 7811 12480 7819 12544
rect 7499 11456 7819 12480
rect 7499 11392 7507 11456
rect 7571 11392 7587 11456
rect 7651 11392 7667 11456
rect 7731 11392 7747 11456
rect 7811 11392 7819 11456
rect 7499 11338 7819 11392
rect 7499 11102 7541 11338
rect 7777 11102 7819 11338
rect 7499 10368 7819 11102
rect 7499 10304 7507 10368
rect 7571 10304 7587 10368
rect 7651 10304 7667 10368
rect 7731 10304 7747 10368
rect 7811 10304 7819 10368
rect 7499 9280 7819 10304
rect 7499 9216 7507 9280
rect 7571 9216 7587 9280
rect 7651 9216 7667 9280
rect 7731 9216 7747 9280
rect 7811 9216 7819 9280
rect 7499 8754 7819 9216
rect 7499 8518 7541 8754
rect 7777 8518 7819 8754
rect 7499 8192 7819 8518
rect 7499 8128 7507 8192
rect 7571 8128 7587 8192
rect 7651 8128 7667 8192
rect 7731 8128 7747 8192
rect 7811 8128 7819 8192
rect 7499 7104 7819 8128
rect 7499 7040 7507 7104
rect 7571 7040 7587 7104
rect 7651 7040 7667 7104
rect 7731 7040 7747 7104
rect 7811 7040 7819 7104
rect 7499 6170 7819 7040
rect 7499 6016 7541 6170
rect 7777 6016 7819 6170
rect 7499 5952 7507 6016
rect 7811 5952 7819 6016
rect 7499 5934 7541 5952
rect 7777 5934 7819 5952
rect 7499 4928 7819 5934
rect 7499 4864 7507 4928
rect 7571 4864 7587 4928
rect 7651 4864 7667 4928
rect 7731 4864 7747 4928
rect 7811 4864 7819 4928
rect 7499 3840 7819 4864
rect 7499 3776 7507 3840
rect 7571 3776 7587 3840
rect 7651 3776 7667 3840
rect 7731 3776 7747 3840
rect 7811 3776 7819 3840
rect 7499 3586 7819 3776
rect 7499 3350 7541 3586
rect 7777 3350 7819 3586
rect 7499 2752 7819 3350
rect 7499 2688 7507 2752
rect 7571 2688 7587 2752
rect 7651 2688 7667 2752
rect 7731 2688 7747 2752
rect 7811 2688 7819 2752
rect 7499 2128 7819 2688
rect 8159 12000 8479 12560
rect 8159 11936 8167 12000
rect 8231 11998 8247 12000
rect 8311 11998 8327 12000
rect 8391 11998 8407 12000
rect 8471 11936 8479 12000
rect 8159 11762 8201 11936
rect 8437 11762 8479 11936
rect 8159 10912 8479 11762
rect 8159 10848 8167 10912
rect 8231 10848 8247 10912
rect 8311 10848 8327 10912
rect 8391 10848 8407 10912
rect 8471 10848 8479 10912
rect 8159 9824 8479 10848
rect 8159 9760 8167 9824
rect 8231 9760 8247 9824
rect 8311 9760 8327 9824
rect 8391 9760 8407 9824
rect 8471 9760 8479 9824
rect 8159 9414 8479 9760
rect 8159 9178 8201 9414
rect 8437 9178 8479 9414
rect 8159 8736 8479 9178
rect 8159 8672 8167 8736
rect 8231 8672 8247 8736
rect 8311 8672 8327 8736
rect 8391 8672 8407 8736
rect 8471 8672 8479 8736
rect 8159 7648 8479 8672
rect 8159 7584 8167 7648
rect 8231 7584 8247 7648
rect 8311 7584 8327 7648
rect 8391 7584 8407 7648
rect 8471 7584 8479 7648
rect 8159 6830 8479 7584
rect 8159 6594 8201 6830
rect 8437 6594 8479 6830
rect 8159 6560 8479 6594
rect 8159 6496 8167 6560
rect 8231 6496 8247 6560
rect 8311 6496 8327 6560
rect 8391 6496 8407 6560
rect 8471 6496 8479 6560
rect 8159 5472 8479 6496
rect 8159 5408 8167 5472
rect 8231 5408 8247 5472
rect 8311 5408 8327 5472
rect 8391 5408 8407 5472
rect 8471 5408 8479 5472
rect 8159 4384 8479 5408
rect 8159 4320 8167 4384
rect 8231 4320 8247 4384
rect 8311 4320 8327 4384
rect 8391 4320 8407 4384
rect 8471 4320 8479 4384
rect 8159 4246 8479 4320
rect 8159 4010 8201 4246
rect 8437 4010 8479 4246
rect 8159 3296 8479 4010
rect 8159 3232 8167 3296
rect 8231 3232 8247 3296
rect 8311 3232 8327 3296
rect 8391 3232 8407 3296
rect 8471 3232 8479 3296
rect 8159 2208 8479 3232
rect 8159 2144 8167 2208
rect 8231 2144 8247 2208
rect 8311 2144 8327 2208
rect 8391 2144 8407 2208
rect 8471 2144 8479 2208
rect 8159 2128 8479 2144
rect 10121 12544 10441 12560
rect 10121 12480 10129 12544
rect 10193 12480 10209 12544
rect 10273 12480 10289 12544
rect 10353 12480 10369 12544
rect 10433 12480 10441 12544
rect 10121 11456 10441 12480
rect 10121 11392 10129 11456
rect 10193 11392 10209 11456
rect 10273 11392 10289 11456
rect 10353 11392 10369 11456
rect 10433 11392 10441 11456
rect 10121 11338 10441 11392
rect 10121 11102 10163 11338
rect 10399 11102 10441 11338
rect 10121 10368 10441 11102
rect 10121 10304 10129 10368
rect 10193 10304 10209 10368
rect 10273 10304 10289 10368
rect 10353 10304 10369 10368
rect 10433 10304 10441 10368
rect 10121 9280 10441 10304
rect 10121 9216 10129 9280
rect 10193 9216 10209 9280
rect 10273 9216 10289 9280
rect 10353 9216 10369 9280
rect 10433 9216 10441 9280
rect 10121 8754 10441 9216
rect 10121 8518 10163 8754
rect 10399 8518 10441 8754
rect 10121 8192 10441 8518
rect 10121 8128 10129 8192
rect 10193 8128 10209 8192
rect 10273 8128 10289 8192
rect 10353 8128 10369 8192
rect 10433 8128 10441 8192
rect 10121 7104 10441 8128
rect 10121 7040 10129 7104
rect 10193 7040 10209 7104
rect 10273 7040 10289 7104
rect 10353 7040 10369 7104
rect 10433 7040 10441 7104
rect 10121 6170 10441 7040
rect 10121 6016 10163 6170
rect 10399 6016 10441 6170
rect 10121 5952 10129 6016
rect 10433 5952 10441 6016
rect 10121 5934 10163 5952
rect 10399 5934 10441 5952
rect 10121 4928 10441 5934
rect 10121 4864 10129 4928
rect 10193 4864 10209 4928
rect 10273 4864 10289 4928
rect 10353 4864 10369 4928
rect 10433 4864 10441 4928
rect 10121 3840 10441 4864
rect 10121 3776 10129 3840
rect 10193 3776 10209 3840
rect 10273 3776 10289 3840
rect 10353 3776 10369 3840
rect 10433 3776 10441 3840
rect 10121 3586 10441 3776
rect 10121 3350 10163 3586
rect 10399 3350 10441 3586
rect 10121 2752 10441 3350
rect 10121 2688 10129 2752
rect 10193 2688 10209 2752
rect 10273 2688 10289 2752
rect 10353 2688 10369 2752
rect 10433 2688 10441 2752
rect 10121 2128 10441 2688
rect 10781 12000 11101 12560
rect 10781 11936 10789 12000
rect 10853 11998 10869 12000
rect 10933 11998 10949 12000
rect 11013 11998 11029 12000
rect 11093 11936 11101 12000
rect 10781 11762 10823 11936
rect 11059 11762 11101 11936
rect 10781 10912 11101 11762
rect 10781 10848 10789 10912
rect 10853 10848 10869 10912
rect 10933 10848 10949 10912
rect 11013 10848 11029 10912
rect 11093 10848 11101 10912
rect 10781 9824 11101 10848
rect 10781 9760 10789 9824
rect 10853 9760 10869 9824
rect 10933 9760 10949 9824
rect 11013 9760 11029 9824
rect 11093 9760 11101 9824
rect 10781 9414 11101 9760
rect 10781 9178 10823 9414
rect 11059 9178 11101 9414
rect 10781 8736 11101 9178
rect 10781 8672 10789 8736
rect 10853 8672 10869 8736
rect 10933 8672 10949 8736
rect 11013 8672 11029 8736
rect 11093 8672 11101 8736
rect 10781 7648 11101 8672
rect 10781 7584 10789 7648
rect 10853 7584 10869 7648
rect 10933 7584 10949 7648
rect 11013 7584 11029 7648
rect 11093 7584 11101 7648
rect 10781 6830 11101 7584
rect 10781 6594 10823 6830
rect 11059 6594 11101 6830
rect 10781 6560 11101 6594
rect 10781 6496 10789 6560
rect 10853 6496 10869 6560
rect 10933 6496 10949 6560
rect 11013 6496 11029 6560
rect 11093 6496 11101 6560
rect 10781 5472 11101 6496
rect 10781 5408 10789 5472
rect 10853 5408 10869 5472
rect 10933 5408 10949 5472
rect 11013 5408 11029 5472
rect 11093 5408 11101 5472
rect 10781 4384 11101 5408
rect 10781 4320 10789 4384
rect 10853 4320 10869 4384
rect 10933 4320 10949 4384
rect 11013 4320 11029 4384
rect 11093 4320 11101 4384
rect 10781 4246 11101 4320
rect 10781 4010 10823 4246
rect 11059 4010 11101 4246
rect 10781 3296 11101 4010
rect 10781 3232 10789 3296
rect 10853 3232 10869 3296
rect 10933 3232 10949 3296
rect 11013 3232 11029 3296
rect 11093 3232 11101 3296
rect 10781 2208 11101 3232
rect 10781 2144 10789 2208
rect 10853 2144 10869 2208
rect 10933 2144 10949 2208
rect 11013 2144 11029 2208
rect 11093 2144 11101 2208
rect 10781 2128 11101 2144
<< via4 >>
rect 2297 11102 2533 11338
rect 2297 8518 2533 8754
rect 2297 6016 2533 6170
rect 2297 5952 2327 6016
rect 2327 5952 2343 6016
rect 2343 5952 2407 6016
rect 2407 5952 2423 6016
rect 2423 5952 2487 6016
rect 2487 5952 2503 6016
rect 2503 5952 2533 6016
rect 2297 5934 2533 5952
rect 2297 3350 2533 3586
rect 2957 11936 2987 11998
rect 2987 11936 3003 11998
rect 3003 11936 3067 11998
rect 3067 11936 3083 11998
rect 3083 11936 3147 11998
rect 3147 11936 3163 11998
rect 3163 11936 3193 11998
rect 2957 11762 3193 11936
rect 2957 9178 3193 9414
rect 2957 6594 3193 6830
rect 2957 4010 3193 4246
rect 4919 11102 5155 11338
rect 4919 8518 5155 8754
rect 4919 6016 5155 6170
rect 4919 5952 4949 6016
rect 4949 5952 4965 6016
rect 4965 5952 5029 6016
rect 5029 5952 5045 6016
rect 5045 5952 5109 6016
rect 5109 5952 5125 6016
rect 5125 5952 5155 6016
rect 4919 5934 5155 5952
rect 4919 3350 5155 3586
rect 5579 11936 5609 11998
rect 5609 11936 5625 11998
rect 5625 11936 5689 11998
rect 5689 11936 5705 11998
rect 5705 11936 5769 11998
rect 5769 11936 5785 11998
rect 5785 11936 5815 11998
rect 5579 11762 5815 11936
rect 5579 9178 5815 9414
rect 5579 6594 5815 6830
rect 5579 4010 5815 4246
rect 7541 11102 7777 11338
rect 7541 8518 7777 8754
rect 7541 6016 7777 6170
rect 7541 5952 7571 6016
rect 7571 5952 7587 6016
rect 7587 5952 7651 6016
rect 7651 5952 7667 6016
rect 7667 5952 7731 6016
rect 7731 5952 7747 6016
rect 7747 5952 7777 6016
rect 7541 5934 7777 5952
rect 7541 3350 7777 3586
rect 8201 11936 8231 11998
rect 8231 11936 8247 11998
rect 8247 11936 8311 11998
rect 8311 11936 8327 11998
rect 8327 11936 8391 11998
rect 8391 11936 8407 11998
rect 8407 11936 8437 11998
rect 8201 11762 8437 11936
rect 8201 9178 8437 9414
rect 8201 6594 8437 6830
rect 8201 4010 8437 4246
rect 10163 11102 10399 11338
rect 10163 8518 10399 8754
rect 10163 6016 10399 6170
rect 10163 5952 10193 6016
rect 10193 5952 10209 6016
rect 10209 5952 10273 6016
rect 10273 5952 10289 6016
rect 10289 5952 10353 6016
rect 10353 5952 10369 6016
rect 10369 5952 10399 6016
rect 10163 5934 10399 5952
rect 10163 3350 10399 3586
rect 10823 11936 10853 11998
rect 10853 11936 10869 11998
rect 10869 11936 10933 11998
rect 10933 11936 10949 11998
rect 10949 11936 11013 11998
rect 11013 11936 11029 11998
rect 11029 11936 11059 11998
rect 10823 11762 11059 11936
rect 10823 9178 11059 9414
rect 10823 6594 11059 6830
rect 10823 4010 11059 4246
<< metal5 >>
rect 1056 11998 11640 12040
rect 1056 11762 2957 11998
rect 3193 11762 5579 11998
rect 5815 11762 8201 11998
rect 8437 11762 10823 11998
rect 11059 11762 11640 11998
rect 1056 11720 11640 11762
rect 1056 11338 11640 11380
rect 1056 11102 2297 11338
rect 2533 11102 4919 11338
rect 5155 11102 7541 11338
rect 7777 11102 10163 11338
rect 10399 11102 11640 11338
rect 1056 11060 11640 11102
rect 1056 9414 11640 9456
rect 1056 9178 2957 9414
rect 3193 9178 5579 9414
rect 5815 9178 8201 9414
rect 8437 9178 10823 9414
rect 11059 9178 11640 9414
rect 1056 9136 11640 9178
rect 1056 8754 11640 8796
rect 1056 8518 2297 8754
rect 2533 8518 4919 8754
rect 5155 8518 7541 8754
rect 7777 8518 10163 8754
rect 10399 8518 11640 8754
rect 1056 8476 11640 8518
rect 1056 6830 11640 6872
rect 1056 6594 2957 6830
rect 3193 6594 5579 6830
rect 5815 6594 8201 6830
rect 8437 6594 10823 6830
rect 11059 6594 11640 6830
rect 1056 6552 11640 6594
rect 1056 6170 11640 6212
rect 1056 5934 2297 6170
rect 2533 5934 4919 6170
rect 5155 5934 7541 6170
rect 7777 5934 10163 6170
rect 10399 5934 11640 6170
rect 1056 5892 11640 5934
rect 1056 4246 11640 4288
rect 1056 4010 2957 4246
rect 3193 4010 5579 4246
rect 5815 4010 8201 4246
rect 8437 4010 10823 4246
rect 11059 4010 11640 4246
rect 1056 3968 11640 4010
rect 1056 3586 11640 3628
rect 1056 3350 2297 3586
rect 2533 3350 4919 3586
rect 5155 3350 7541 3586
rect 7777 3350 10163 3586
rect 10399 3350 11640 3586
rect 1056 3308 11640 3350
use sky130_fd_sc_hd__xor2_1  _1_
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2_
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _3_
timestamp 0
transform -1 0 7268 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 0
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_6
timestamp 0
transform 1 0 1656 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_18
timestamp 0
transform 1 0 2760 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_30
timestamp 0
transform 1 0 3864 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_42
timestamp 0
transform 1 0 4968 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_50
timestamp 0
transform 1 0 5704 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_67
timestamp 0
transform 1 0 7268 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_79
timestamp 0
transform 1 0 8372 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_91
timestamp 0
transform 1 0 9476 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_103
timestamp 0
transform 1 0 10580 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_6
timestamp 0
transform 1 0 1656 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_18
timestamp 0
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_26
timestamp 0
transform 1 0 3496 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_105
timestamp 0
transform 1 0 10764 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_57
timestamp 0
transform 1 0 6348 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_69
timestamp 0
transform 1 0 7452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_81
timestamp 0
transform 1 0 8556 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output3
timestamp 0
transform 1 0 10948 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output4
timestamp 0
transform 1 0 10948 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_19
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 0
transform -1 0 11592 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_20
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 0
transform -1 0 11592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_21
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 0
transform -1 0 11592 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_22
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 0
transform -1 0 11592 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_23
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 0
transform -1 0 11592 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_24
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 0
transform -1 0 11592 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_25
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 0
transform -1 0 11592 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_26
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 0
transform -1 0 11592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_27
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 0
transform -1 0 11592 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_28
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 0
transform -1 0 11592 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_29
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 0
transform -1 0 11592 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_30
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 0
transform -1 0 11592 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_31
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 0
transform -1 0 11592 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_32
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 0
transform -1 0 11592 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_33
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 0
transform -1 0 11592 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_34
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 0
transform -1 0 11592 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_35
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 0
transform -1 0 11592 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_36
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 0
transform -1 0 11592 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_37
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 0
transform -1 0 11592 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_38
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_39
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_40
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_41
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_42
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_43
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_44
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_45
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_46
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_47
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_48
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_49
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_50
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_51
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_52
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_53
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_54
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_55
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_56
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_57
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_58
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_59
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_60
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_61
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_62
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_63
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_64
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_65
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_66
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_67
timestamp 0
transform 1 0 6256 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_68
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
<< labels >>
rlabel metal1 s 6348 11968 6348 11968 4 VGND
rlabel metal1 s 6348 12512 6348 12512 4 VPWR
rlabel metal1 s 6555 7514 6555 7514 4 _0_
rlabel metal3 s 1050 6868 1050 6868 4 in1
rlabel metal3 s 0 7488 800 7608 4 in4
port 4 nsew
rlabel metal1 s 6026 7344 6026 7344 4 net1
rlabel metal1 s 3726 7378 3726 7378 4 net2
rlabel metal2 s 7222 7684 7222 7684 4 net3
rlabel metal1 s 8970 7310 8970 7310 4 net4
rlabel metal1 s 11224 7718 11224 7718 4 out2
rlabel metal3 s 11600 6868 11600 6868 4 out3
flabel metal5 s 1056 11720 11640 12040 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 9136 11640 9456 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6552 11640 6872 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 3968 11640 4288 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 10781 2128 11101 12560 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 8159 2128 8479 12560 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5537 2128 5857 12560 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 2915 2128 3235 12560 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 11060 11640 11380 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 8476 11640 8796 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5892 11640 6212 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 3308 11640 3628 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 10121 2128 10441 12560 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 7499 2128 7819 12560 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4877 2128 5197 12560 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 2255 2128 2575 12560 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 0 6808 800 6928 0 FreeSans 600 0 0 0 in1
port 3 nsew
flabel metal3 s 400 7548 400 7548 0 FreeSans 600 0 0 0 in4
flabel metal3 s 11901 7488 12701 7608 0 FreeSans 600 0 0 0 out2
port 5 nsew
flabel metal3 s 11901 6808 12701 6928 0 FreeSans 600 0 0 0 out3
port 6 nsew
<< properties >>
string FIXED_BBOX 0 0 12701 14845
<< end >>
