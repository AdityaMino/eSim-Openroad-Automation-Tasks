magic
tech sky130A
magscale 1 2
timestamp 1750272434
<< nwell >>
rect 1066 2159 11630 12550
<< obsli1 >>
rect 1104 2159 11592 12529
<< obsm1 >>
rect 842 2128 11592 12560
<< obsm2 >>
rect 846 2139 11298 12549
<< metal3 >>
rect 0 7488 800 7608
rect 11901 7488 12701 7608
rect 0 6808 800 6928
rect 11901 6808 12701 6928
<< obsm3 >>
rect 798 7688 11901 12545
rect 880 7408 11821 7688
rect 798 7008 11901 7408
rect 880 6728 11821 7008
rect 798 2143 11901 6728
<< metal4 >>
rect 2255 2128 2575 12560
rect 2915 2128 3235 12560
rect 4877 2128 5197 12560
rect 5537 2128 5857 12560
rect 7499 2128 7819 12560
rect 8159 2128 8479 12560
rect 10121 2128 10441 12560
rect 10781 2128 11101 12560
<< metal5 >>
rect 1056 11720 11640 12040
rect 1056 11060 11640 11380
rect 1056 9136 11640 9456
rect 1056 8476 11640 8796
rect 1056 6552 11640 6872
rect 1056 5892 11640 6212
rect 1056 3968 11640 4288
rect 1056 3308 11640 3628
<< labels >>
rlabel metal4 s 2915 2128 3235 12560 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 5537 2128 5857 12560 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 8159 2128 8479 12560 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 10781 2128 11101 12560 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 3968 11640 4288 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6552 11640 6872 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9136 11640 9456 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 11720 11640 12040 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 2255 2128 2575 12560 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 4877 2128 5197 12560 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7499 2128 7819 12560 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 10121 2128 10441 12560 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 3308 11640 3628 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5892 11640 6212 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8476 11640 8796 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11060 11640 11380 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 6808 800 6928 6 in1
port 3 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 in4
port 4 nsew signal input
rlabel metal3 s 11901 7488 12701 7608 6 out2
port 5 nsew signal output
rlabel metal3 s 11901 6808 12701 6928 6 out3
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 12701 14845
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 159626
string GDS_FILE /openlane/designs/halfadder/runs/RUN_2025.06.18_18.46.26/results/signoff/halfadder.magic.gds
string GDS_START 42988
<< end >>

